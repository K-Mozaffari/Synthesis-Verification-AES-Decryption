
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_aes_dec_KEY_SIZE2 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_aes_dec_KEY_SIZE2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_aes_dec_KEY_SIZE2.all;

entity key_expansion is

   port( KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, CLK_I, RESET_I
         , CE_I : in std_logic;  DONE_O : out std_logic;  GET_KEY_I : in 
         std_logic;  KEY_NUMB_I : in std_logic_vector (5 downto 0);  KEY_EXP_O 
         : out std_logic_vector (31 downto 0));

end key_expansion;

architecture SYN_Behavioral of key_expansion is

   component IVI
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EO
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EN
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ND3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO7
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EON1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component NR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component IVDA
      port( A : in std_logic;  Y, Z : out std_logic);
   end component;
   
   component EOI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AN2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2P
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component B2I
      port( A : in std_logic;  Z1, Z2 : out std_logic);
   end component;
   
   component NR3P
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO1P
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component IVDAP
      port( A : in std_logic;  Y, Z : out std_logic);
   end component;
   
   component B3IP
      port( A : in std_logic;  Z1, Z2 : out std_logic);
   end component;
   
   component AN3P
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ENI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2P
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FD1
      port( D, CP : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal v_KEY32_IN_31_port, v_KEY32_IN_30_port, v_KEY32_IN_29_port, 
      v_KEY32_IN_28_port, v_KEY32_IN_27_port, v_KEY32_IN_26_port, 
      v_KEY32_IN_25_port, v_KEY32_IN_24_port, v_KEY32_IN_23_port, 
      v_KEY32_IN_22_port, v_KEY32_IN_21_port, v_KEY32_IN_20_port, 
      v_KEY32_IN_19_port, v_KEY32_IN_18_port, v_KEY32_IN_17_port, 
      v_KEY32_IN_16_port, v_KEY32_IN_15_port, v_KEY32_IN_14_port, 
      v_KEY32_IN_13_port, v_KEY32_IN_12_port, v_KEY32_IN_11_port, 
      v_KEY32_IN_10_port, v_KEY32_IN_9_port, v_KEY32_IN_8_port, 
      v_KEY32_IN_7_port, v_KEY32_IN_6_port, v_KEY32_IN_5_port, 
      v_KEY32_IN_4_port, v_KEY32_IN_3_port, v_KEY32_IN_2_port, 
      v_KEY32_IN_1_port, v_KEY32_IN_0_port, v_CALCULATION_CNTR_7_port, 
      v_CALCULATION_CNTR_6_port, v_CALCULATION_CNTR_5_port, 
      v_CALCULATION_CNTR_4_port, v_CALCULATION_CNTR_3_port, 
      v_CALCULATION_CNTR_2_port, v_CALCULATION_CNTR_1_port, 
      v_CALCULATION_CNTR_0_port, i_SRAM_ADDR_WR0_5_port, i_SRAM_ADDR_WR0_4_port
      , i_SRAM_ADDR_WR0_3_port, i_SRAM_ADDR_WR0_2_port, i_SRAM_ADDR_WR0_1_port,
      i_SRAM_ADDR_WR0_0_port, v_KEY_COL_OUT0_31_port, v_KEY_COL_OUT0_30_port, 
      v_KEY_COL_OUT0_29_port, v_KEY_COL_OUT0_28_port, v_KEY_COL_OUT0_27_port, 
      v_KEY_COL_OUT0_26_port, v_KEY_COL_OUT0_25_port, v_KEY_COL_OUT0_24_port, 
      v_KEY_COL_OUT0_23_port, v_KEY_COL_OUT0_22_port, v_KEY_COL_OUT0_21_port, 
      v_KEY_COL_OUT0_20_port, v_KEY_COL_OUT0_19_port, v_KEY_COL_OUT0_18_port, 
      v_KEY_COL_OUT0_17_port, v_KEY_COL_OUT0_16_port, v_KEY_COL_OUT0_15_port, 
      v_KEY_COL_OUT0_14_port, v_KEY_COL_OUT0_13_port, v_KEY_COL_OUT0_12_port, 
      v_KEY_COL_OUT0_11_port, v_KEY_COL_OUT0_10_port, v_KEY_COL_OUT0_9_port, 
      v_KEY_COL_OUT0_8_port, i_INTERN_ADDR_RD0_5_port, i_INTERN_ADDR_RD0_4_port
      , i_INTERN_ADDR_RD0_3_port, i_INTERN_ADDR_RD0_2_port, 
      i_INTERN_ADDR_RD0_1_port, i_INTERN_ADDR_RD0_0_port, v_TEMP_VECTOR_31_port
      , v_TEMP_VECTOR_30_port, v_TEMP_VECTOR_29_port, v_TEMP_VECTOR_28_port, 
      v_TEMP_VECTOR_27_port, v_TEMP_VECTOR_26_port, v_TEMP_VECTOR_25_port, 
      v_TEMP_VECTOR_24_port, v_TEMP_VECTOR_23_port, v_TEMP_VECTOR_22_port, 
      v_TEMP_VECTOR_21_port, v_TEMP_VECTOR_20_port, v_TEMP_VECTOR_19_port, 
      v_TEMP_VECTOR_18_port, v_TEMP_VECTOR_17_port, v_TEMP_VECTOR_16_port, 
      v_TEMP_VECTOR_15_port, v_TEMP_VECTOR_14_port, v_TEMP_VECTOR_13_port, 
      v_TEMP_VECTOR_12_port, v_TEMP_VECTOR_11_port, v_TEMP_VECTOR_10_port, 
      v_TEMP_VECTOR_9_port, v_TEMP_VECTOR_8_port, v_TEMP_VECTOR_7_port, 
      v_TEMP_VECTOR_6_port, v_TEMP_VECTOR_5_port, v_TEMP_VECTOR_4_port, 
      v_TEMP_VECTOR_3_port, v_TEMP_VECTOR_2_port, v_TEMP_VECTOR_1_port, 
      v_TEMP_VECTOR_0_port, v_SUB_WORD_7_port, N1748, N1749, N1750, N1751, 
      N1752, N1753, N1754, n13, n15, n16, n17, n18, n19, n20, n21, n24, n25, 
      n26, n27, n29, n30, n31, n32, n34, n35, n36, n37, n39, n40, n41, n42, n44
      , n45, n46, n47, n49, n50, n51, n52, n54, n55, n56, n57, n58, n60, n61, 
      n62, n64, n65, n66, n67, n68, n70, n73, n74, n75, n76, n77, n78, n79, n80
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n164, n165, n166, n167, n168, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n183, n184, n185, n186, n187, n189, n190, 
      n191, n192, n193, n194, n195, n197, n199, n200, n201, n202, n203, n205, 
      n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218, n219, 
      n220, n222, n223, n225, n226, n227, n228, n229, n230, n231, n232, n236, 
      n237, n239, n245, n246, n249, n250, n253, n257, n258, n259, n260, n262, 
      n268, n270, n272, n275, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n289, n291, n292, n293, n295, n296, n298, n299, n300, 
      n301, n302, n303, n304, n305, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n359, n360, 
      n361, n362, n371, n372, n373, n374, n383, n384, n385, n386, n395, n396, 
      n397, n398, n399, n400, n401, n402, n411, n412, n413, n414, n423, n424, 
      n425, n426, n435, n436, n437, n438, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
      n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n843, n844, n845, 
      n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, 
      n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, 
      n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, 
      n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, 
      n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, 
      n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, 
      n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
      n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
      n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1149, n1150, n1151, n1152, n1153, n1154, n1155, 
      n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, 
      n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, 
      n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, 
      n1186, n1187, n1188, n1189, n1190, n1191, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
      n1450, n1451, n1452, n1453, n1455, n1456, n1457, n1458, n1459, n1460, 
      n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
      n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
      n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, 
      n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1499, n1500, n1501, 
      n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, 
      n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
      n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
      n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
      n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, 
      n1624, n1625, n1626, n1627, n1628, n1629, n1631, n1632, n1633, n1634, 
      n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, 
      n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
      n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, 
      n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748_port, n1749_port, n1750_port, n1751_port, n1752_port, 
      n1753_port, n1754_port, n1755, n1756, n1757, n1758, n1759, n1760, n1761, 
      n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
      n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, 
      n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1792, n1793, 
      n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1824, n1825, n1826, n1827, n1828, n1829, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1840, n1843, n1844, n1846, n1847, n1849, 
      n1850, n1851, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, 
      n1861, n1863, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, 
      n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1884, 
      n1886, n1888, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1898, 
      n1899, n1900, n1901, n1902, n1905, n1908, n1911, n1912, n1913, n1914, 
      n1915, n1916, n1917, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1944, n1945, n1946, n1948, n1949, n1950, n1951, 
      n1952, n1956, n1957, n1958, n1961, n1962, n1963, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1975, n1977, n1979, n1980, 
      n1981, n1982, n1983, n1984, n1987, n1988, n1990, n1991, n1993, n1994, 
      n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2007, 
      n2008, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2028, n2029, 
      n2030, n2031, n2032, n2034, n2036, n2038, n2039, n2040, n2041, n2042, 
      n2044, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
      n2056, n2057, n2058, n2060, n2061, n2062, n2063, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2082, n2083, n2084, n2086, n2087, n2088, n2089, 
      n2090, n2091, n2093, n2094, n2096, n2097, n2098, n2099, n2100, n2101, 
      n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, 
      n2134, n2135, n2137, n2138, n2139, n2141, n2142, n2143, n2144, n2145, 
      n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, 
      n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
      n2167, n2170, n2171, n2172, n2173, n2175, n2176, n2177, n2178, n2179, 
      n2180, n2181, n2182, n2184, n2185, n2186, n2187, n2188, n2190, n2191, 
      n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2201, n2202, 
      n2203, n2204, n2205, n2207, n2208, n2209, n2210, n2211, n2212, n2213, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, 
      n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2235, 
      n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
      n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
      n2257, n2258, n2259, n2260, n2261, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2289, n2291, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
      n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
      n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
      n2462, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2475, n2476, n2477, n2478, n2479, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2491, n2492, n2493, n2494, n2495, n2496, n2497, 
      n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, 
      n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
      n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, 
      n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, 
      n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, 
      n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, 
      n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, 
      n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, 
      n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
      n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, 
      n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, 
      n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, 
      n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
      n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
      n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, 
      n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, 
      n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, 
      n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, 
      n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, 
      n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
      n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, 
      n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
      n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
      n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, 
      n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, 
      n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, 
      n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, 
      n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, 
      n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, 
      n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, 
      n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, 
      n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
      n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, 
      n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, 
      n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, 
      n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, 
      n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, 
      n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, 
      n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, 
      n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, 
      n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, 
      n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, 
      n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, 
      n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, 
      n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, 
      n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
      n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
      n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, 
      n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
      n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, 
      n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
      n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, 
      n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, 
      n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, 
      n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, 
      n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, 
      n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, 
      n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
      n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, 
      n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
      n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, 
      n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, 
      n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, 
      n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, 
      n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, 
      n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, 
      n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, 
      n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, 
      n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, 
      n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, 
      n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, 
      n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, 
      n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, 
      n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, 
      n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, 
      n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, 
      n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, 
      n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, 
      n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, 
      n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, 
      n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, 
      n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, 
      n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, 
      n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, 
      n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, 
      n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, 
      n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, 
      n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, 
      n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, 
      n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, 
      n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, 
      n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, 
      n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, 
      n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, 
      n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, 
      n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, 
      n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, 
      n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, 
      n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, 
      n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, 
      n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, 
      n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, 
      n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, 
      n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, 
      n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, 
      n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
      n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, 
      n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, 
      n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, 
      n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, 
      n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, 
      n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, 
      n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, 
      n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, 
      n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, 
      n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, 
      n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, 
      n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, 
      n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, 
      n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, 
      n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, 
      n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, 
      n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, 
      n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, 
      n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, 
      n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, 
      n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, 
      n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, 
      n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, 
      n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, 
      n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, 
      n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, 
      n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, 
      n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, 
      n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, 
      n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, 
      n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, 
      n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, 
      n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, 
      n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, 
      n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, 
      n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, 
      n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, 
      n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, 
      n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, 
      n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, 
      n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, 
      n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, 
      n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, 
      n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, 
      n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, 
      n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
      n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
      n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
      n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
      n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, 
      n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
      n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, 
      n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, 
      n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, 
      n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, 
      n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, 
      n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, 
      n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, 
      n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
      n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, 
      n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, 
      n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, 
      n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, 
      n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, 
      n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, 
      n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, 
      n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
      n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4544, n4545, n4546, n4547, n4548, n4549, 
      n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, 
      n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, 
      n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, 
      n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, 
      n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, 
      n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, 
      n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, 
      n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, 
      n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, 
      n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, 
      n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, 
      n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, 
      n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, 
      n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, 
      n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, 
      n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, 
      n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, 
      n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, 
      n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, 
      n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, 
      n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, 
      n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, 
      n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, 
      n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, 
      n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, 
      n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, 
      n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, 
      n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, 
      n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, 
      n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, 
      n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, 
      n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, 
      n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, 
      n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, 
      n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, 
      n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, 
      n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, 
      n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, 
      n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, 
      n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, 
      n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, 
      n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, 
      n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, 
      n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, 
      n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, 
      n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, 
      n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, 
      n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, 
      n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, 
      n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, 
      n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, 
      n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, 
      n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, 
      n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, 
      n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, 
      n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, 
      n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, 
      n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, 
      n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, 
      n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, 
      n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, 
      n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, 
      n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, 
      n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, 
      n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, 
      n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, 
      n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, 
      n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, 
      n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, 
      n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, 
      n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, 
      n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, 
      n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, 
      n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, 
      n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, 
      n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
      n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, 
      n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, 
      n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
      n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, 
      n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, 
      n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, 
      n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, 
      n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, 
      n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, 
      n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, 
      n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, 
      n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, 
      n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, 
      n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, 
      n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, 
      n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
      n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, 
      n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, 
      n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, 
      n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, 
      n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, 
      n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, 
      n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, 
      n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, 
      n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, 
      n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, 
      n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, 
      n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, 
      n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, 
      n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, 
      n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, 
      n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, 
      n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, 
      n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, 
      n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, 
      n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, 
      n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, 
      n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, 
      n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, 
      n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, 
      n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, 
      n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, 
      n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, 
      n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, 
      n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, 
      n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, 
      n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, 
      n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, 
      n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, 
      n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, 
      n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, 
      n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, 
      n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, 
      n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, 
      n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, 
      n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, 
      n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, 
      n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, 
      n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, 
      n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, 
      n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, 
      n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, 
      n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, 
      n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, 
      n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, 
      n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, 
      n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, 
      n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, 
      n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, 
      n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, 
      n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, 
      n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, 
      n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, 
      n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, 
      n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, 
      n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, 
      n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, 
      n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, 
      n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, 
      n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, 
      n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, 
      n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, 
      n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, 
      n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, 
      n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, 
      n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, 
      n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, 
      n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, 
      n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, 
      n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, 
      n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, 
      n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, 
      n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, 
      n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, 
      n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, 
      n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, 
      n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, 
      n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, 
      n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, 
      n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, 
      n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, 
      n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, 
      n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, 
      n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, 
      n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, 
      n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, 
      n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, 
      n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, 
      n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, 
      n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, 
      n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, 
      n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, 
      n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, 
      n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, 
      n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, 
      n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, 
      n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, 
      n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, 
      n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, 
      n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, 
      n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, 
      n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, 
      n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, 
      n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, 
      n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, 
      n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, 
      n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, 
      n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, 
      n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, 
      n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, 
      n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, 
      n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, 
      n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, 
      n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, 
      n6651, n6652, n6653, n6654, n6655, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6748, n6749, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
      n12, n14, n22, n23, n28, n33, n38, n43, n48, n53, n59, n63, n69, n71, n72
      , n81, n109, n122, n150, n163, n169, n170, n171, n181, n182, n188, n196, 
      n198, n204, n206, n213, n221, n224, n233, n234, n235, n238, n240, n241, 
      n242, n243, n244, n247, n248, n251, n252, n254, n255, n256, n261, n263, 
      n264, n265, n266, n267, n269, n271, n273, n274, n276, n288, n290, n294, 
      n297, n306, n317, n327, n339, n351, n352, n353, n354, n355, n356, n357, 
      n358, n363, n364, n365, n366, n367, n368, n369, n370, n375, n376, n377, 
      n378, n379, n380, n381, n382, n387, n388, n389, n390, n391, n392, n393, 
      n394, n403, n404, n405, n406, n407, n408, n409, n410, n415, n416, n417, 
      n418, n419, n420, n421, n422, n427, n428, n429, n430, n431, n432, n433, 
      n434, n439, n440, n441, n442, n443, n444, n445, n446, n447, n491, n535, 
      n579, n623, n667, n754, n798, n842, n929, n973, n1017, n1104, n1148, 
      n1192, n1279, n1323, n1367, n1454, n1498, n1542, n1586, n1630, n1674, 
      n1718, n1790, n1791, n1830, n1831, n1841, n1842, n1845, n1848, n1852, 
      n1862, n1864, n1865, n1883, n1885, n1887, n1889, n1897, n1903, n1904, 
      n1906, n1907, n1909, n1910, n1918, n1919, n1920, n1921, n1932, n1943, 
      n1947, n1953, n1954, n1955, n1959, n1960, n1964, n1974, n1976, n1978, 
      n1985, n1986, n1989, n1992, n2004, n2005, n2006, n2009, n2027, n2033, 
      n2035, n2037, n2043, n2045, n2055, n2059, n2064, n2081, n2085, n2092, 
      n2095, n2111, n2125, n2136, n2140, n2166, n2168, n2169, n2174, n2183, 
      n2189, n2200, n2206, n2214, n2234, n2256, n2262, n2279, n2287, n2288, 
      n2290, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
      n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, 
      n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
      n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, 
      n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
      n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, 
      n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
      n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
      n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
      n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2461, n2463, n2473, n2474, n2480, n2481, n2490, n4542, n4543, n6650, 
      n6656, n6657, n6658, n6716, n6717, n6718, n6719, n6720, n6721, n6722, 
      n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, 
      n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, 
      n6743, n6744, n6745, n6746, n6747, n6750, n6751, n6752, n6753, n6754, 
      n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, 
      n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, 
      n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, 
      n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, 
      n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, 
      n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, 
      n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, 
      n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, 
      n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, 
      n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, 
      n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, 
      n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, 
      n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, 
      n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, 
      n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, 
      n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, 
      n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, 
      n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, 
      n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, 
      n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, 
      n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, 
      n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, 
      n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, 
      n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, 
      n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, 
      n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, 
      n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, 
      n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, 
      n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, 
      n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, 
      n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, 
      n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, 
      n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, 
      n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, 
      n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, 
      n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, 
      n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, 
      n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, 
      n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, 
      n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, 
      n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, 
      n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, 
      n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, 
      n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, 
      n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, 
      n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, 
      n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, 
      n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, 
      n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, 
      n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, 
      n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, 
      n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, 
      n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, 
      n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, 
      n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, 
      n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, 
      n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, 
      n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, 
      n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, 
      n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, 
      n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, 
      n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, 
      n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, 
      n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, 
      n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, 
      n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, 
      n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, 
      n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, 
      n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, 
      n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, 
      n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, 
      n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, 
      n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, 
      n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, 
      n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, 
      n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, 
      n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, 
      n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, 
      n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, 
      n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, 
      n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, 
      n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, 
      n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, 
      n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, 
      n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, 
      n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, 
      n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, 
      n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, 
      n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, 
      n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, 
      n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, 
      n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, 
      n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, 
      n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, 
      n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, 
      n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, 
      n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, 
      n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, 
      n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, 
      n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, 
      n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, 
      n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, 
      n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, 
      n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, 
      n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, 
      n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, 
      n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, 
      n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, 
      n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, 
      n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, 
      n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, 
      n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, 
      n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, 
      n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, 
      n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, 
      n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, 
      n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, 
      n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, 
      n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, 
      n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, 
      n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, 
      n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, 
      n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, 
      n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, 
      n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, 
      n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, 
      n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, 
      n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, 
      n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, 
      n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, 
      n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, 
      n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, 
      n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, 
      n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, 
      n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, 
      n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, 
      n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, 
      n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, 
      n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, 
      n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, 
      n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, 
      n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, 
      n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, 
      n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, 
      n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, 
      n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, 
      n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, 
      n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, 
      n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, 
      n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, 
      n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, 
      n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, 
      n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, 
      n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, 
      n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n_1000, n_1001, 
      n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, 
      n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, 
      n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, 
      n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, 
      n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, 
      n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, 
      n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, 
      n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, 
      n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, 
      n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, 
      n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, 
      n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, 
      n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, 
      n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, 
      n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, 
      n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, 
      n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, 
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, 
      n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, 
      n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, 
      n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, 
      n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, 
      n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, 
      n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, 
      n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, 
      n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, 
      n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, 
      n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, 
      n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, 
      n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, 
      n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, 
      n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, 
      n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, 
      n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, 
      n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, 
      n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, 
      n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, 
      n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, 
      n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, 
      n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, 
      n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, 
      n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, 
      n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, 
      n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, 
      n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, 
      n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, 
      n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, 
      n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, 
      n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, 
      n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, 
      n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, 
      n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, 
      n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, 
      n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, 
      n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, 
      n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, 
      n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, 
      n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, 
      n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, 
      n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, 
      n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, 
      n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, 
      n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, 
      n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, 
      n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, 
      n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, 
      n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, 
      n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, 
      n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, 
      n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, 
      n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, 
      n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, 
      n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, 
      n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, 
      n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, 
      n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, 
      n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, 
      n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, 
      n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, 
      n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, 
      n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, 
      n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, 
      n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, 
      n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, 
      n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, 
      n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, 
      n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, 
      n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, 
      n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, 
      n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, 
      n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, 
      n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, 
      n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, 
      n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, 
      n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, 
      n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, 
      n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, 
      n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, 
      n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, 
      n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, 
      n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, 
      n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, 
      n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, 
      n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, 
      n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, 
      n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, 
      n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, 
      n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, 
      n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, 
      n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, 
      n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, 
      n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, 
      n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, 
      n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, 
      n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, 
      n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, 
      n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, 
      n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, 
      n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, 
      n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, 
      n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, 
      n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, 
      n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, 
      n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, 
      n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, 
      n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, 
      n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, 
      n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, 
      n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, 
      n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, 
      n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, 
      n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, 
      n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, 
      n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, 
      n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, 
      n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, 
      n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, 
      n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, 
      n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, 
      n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, 
      n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, 
      n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, 
      n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, 
      n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, 
      n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, 
      n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, 
      n_3135, n_3136 : std_logic;

begin
   
   i_BYTE_CNTR4_reg_0_inst : FD1 port map( D => n6749, CP => CLK_I, Q => n288, 
                           QN => n2487);
   i_BYTE_CNTR4_reg_1_inst : FD1 port map( D => n6748, CP => CLK_I, Q => n358, 
                           QN => n2488);
   FF_VALID_KEY_reg : FD1 port map( D => n4589, CP => CLK_I, Q => n_1000, QN =>
                           n4548);
   v_KEY32_IN_reg_31_inst : FD1 port map( D => n8188, CP => CLK_I, Q => 
                           v_KEY32_IN_31_port, QN => n_1001);
   v_KEY32_IN_reg_30_inst : FD1 port map( D => n8187, CP => CLK_I, Q => 
                           v_KEY32_IN_30_port, QN => n_1002);
   v_KEY32_IN_reg_29_inst : FD1 port map( D => n8186, CP => CLK_I, Q => 
                           v_KEY32_IN_29_port, QN => n_1003);
   v_KEY32_IN_reg_28_inst : FD1 port map( D => n8185, CP => CLK_I, Q => 
                           v_KEY32_IN_28_port, QN => n_1004);
   v_KEY32_IN_reg_27_inst : FD1 port map( D => n8184, CP => CLK_I, Q => 
                           v_KEY32_IN_27_port, QN => n_1005);
   v_KEY32_IN_reg_26_inst : FD1 port map( D => n8183, CP => CLK_I, Q => 
                           v_KEY32_IN_26_port, QN => n_1006);
   v_KEY32_IN_reg_25_inst : FD1 port map( D => n8182, CP => CLK_I, Q => 
                           v_KEY32_IN_25_port, QN => n_1007);
   v_KEY32_IN_reg_24_inst : FD1 port map( D => n8181, CP => CLK_I, Q => 
                           v_KEY32_IN_24_port, QN => n_1008);
   v_KEY32_IN_reg_23_inst : FD1 port map( D => n8205, CP => CLK_I, Q => 
                           v_KEY32_IN_23_port, QN => n_1009);
   v_KEY32_IN_reg_22_inst : FD1 port map( D => n8204, CP => CLK_I, Q => 
                           v_KEY32_IN_22_port, QN => n_1010);
   v_KEY32_IN_reg_21_inst : FD1 port map( D => n8203, CP => CLK_I, Q => 
                           v_KEY32_IN_21_port, QN => n_1011);
   v_KEY32_IN_reg_20_inst : FD1 port map( D => n8202, CP => CLK_I, Q => 
                           v_KEY32_IN_20_port, QN => n_1012);
   v_KEY32_IN_reg_19_inst : FD1 port map( D => n8201, CP => CLK_I, Q => 
                           v_KEY32_IN_19_port, QN => n_1013);
   v_KEY32_IN_reg_18_inst : FD1 port map( D => n8200, CP => CLK_I, Q => 
                           v_KEY32_IN_18_port, QN => n_1014);
   v_KEY32_IN_reg_17_inst : FD1 port map( D => n8199, CP => CLK_I, Q => 
                           v_KEY32_IN_17_port, QN => n_1015);
   v_KEY32_IN_reg_16_inst : FD1 port map( D => n8198, CP => CLK_I, Q => 
                           v_KEY32_IN_16_port, QN => n_1016);
   v_KEY32_IN_reg_15_inst : FD1 port map( D => n8214, CP => CLK_I, Q => 
                           v_KEY32_IN_15_port, QN => n_1017);
   v_KEY32_IN_reg_14_inst : FD1 port map( D => n8213, CP => CLK_I, Q => 
                           v_KEY32_IN_14_port, QN => n_1018);
   v_KEY32_IN_reg_13_inst : FD1 port map( D => n8212, CP => CLK_I, Q => 
                           v_KEY32_IN_13_port, QN => n_1019);
   v_KEY32_IN_reg_12_inst : FD1 port map( D => n8211, CP => CLK_I, Q => 
                           v_KEY32_IN_12_port, QN => n_1020);
   v_KEY32_IN_reg_11_inst : FD1 port map( D => n8210, CP => CLK_I, Q => 
                           v_KEY32_IN_11_port, QN => n_1021);
   v_KEY32_IN_reg_10_inst : FD1 port map( D => n8209, CP => CLK_I, Q => 
                           v_KEY32_IN_10_port, QN => n_1022);
   v_KEY32_IN_reg_9_inst : FD1 port map( D => n8208, CP => CLK_I, Q => 
                           v_KEY32_IN_9_port, QN => n_1023);
   v_KEY32_IN_reg_8_inst : FD1 port map( D => n8207, CP => CLK_I, Q => 
                           v_KEY32_IN_8_port, QN => n_1024);
   v_KEY32_IN_reg_7_inst : FD1 port map( D => n8197, CP => CLK_I, Q => 
                           v_KEY32_IN_7_port, QN => n_1025);
   v_KEY32_IN_reg_6_inst : FD1 port map( D => n8196, CP => CLK_I, Q => 
                           v_KEY32_IN_6_port, QN => n_1026);
   v_KEY32_IN_reg_5_inst : FD1 port map( D => n8195, CP => CLK_I, Q => 
                           v_KEY32_IN_5_port, QN => n_1027);
   v_KEY32_IN_reg_4_inst : FD1 port map( D => n8194, CP => CLK_I, Q => 
                           v_KEY32_IN_4_port, QN => n_1028);
   v_KEY32_IN_reg_3_inst : FD1 port map( D => n8193, CP => CLK_I, Q => 
                           v_KEY32_IN_3_port, QN => n_1029);
   v_KEY32_IN_reg_2_inst : FD1 port map( D => n8192, CP => CLK_I, Q => 
                           v_KEY32_IN_2_port, QN => n_1030);
   v_KEY32_IN_reg_1_inst : FD1 port map( D => n8191, CP => CLK_I, Q => 
                           v_KEY32_IN_1_port, QN => n_1031);
   v_KEY32_IN_reg_0_inst : FD1 port map( D => n8190, CP => CLK_I, Q => 
                           v_KEY32_IN_0_port, QN => n_1032);
   FF_GET_KEY_reg : FD1 port map( D => GET_KEY_I, CP => CLK_I, Q => n379, QN =>
                           n269);
   v_SUB_WORD_reg_7_inst : FD1 port map( D => n4588, CP => CLK_I, Q => 
                           v_SUB_WORD_7_port, QN => n1960);
   v_SUB_WORD_reg_6_inst : FD1 port map( D => n4587, CP => CLK_I, Q => n_1033, 
                           QN => n1959);
   v_SUB_WORD_reg_5_inst : FD1 port map( D => n4586, CP => CLK_I, Q => n4547, 
                           QN => n1964);
   v_SUB_WORD_reg_4_inst : FD1 port map( D => n4585, CP => CLK_I, Q => n4546, 
                           QN => n1974);
   v_SUB_WORD_reg_3_inst : FD1 port map( D => n4584, CP => CLK_I, Q => n4545, 
                           QN => n1976);
   v_SUB_WORD_reg_2_inst : FD1 port map( D => n4583, CP => CLK_I, Q => n4544, 
                           QN => n1978);
   v_SUB_WORD_reg_1_inst : FD1 port map( D => n4582, CP => CLK_I, Q => n_1034, 
                           QN => n1955);
   v_SUB_WORD_reg_0_inst : FD1 port map( D => n4581, CP => CLK_I, Q => n_1035, 
                           QN => n1954);
   v_CALCULATION_CNTR_reg_0_inst : FD1 port map( D => n6651, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_0_port, QN => n1985);
   i_ROUND_reg_3_inst : FD1 port map( D => n6715, CP => CLK_I, Q => n1921, QN 
                           => n6660);
   START_CALCULATION_reg : FD1 port map( D => n6711, CP => CLK_I, Q => n_1036, 
                           QN => n6659);
   i_ROUND_reg_0_inst : FD1 port map( D => n6714, CP => CLK_I, Q => n290, QN =>
                           n6663);
   i_ROUND_reg_1_inst : FD1 port map( D => n6713, CP => CLK_I, Q => n363, QN =>
                           n6662);
   i_ROUND_reg_2_inst : FD1 port map( D => n6712, CP => CLK_I, Q => n1918, QN 
                           => n6661);
   DONE_O_reg : FD1 port map( D => n6710, CP => CLK_I, Q => DONE_O, QN => n2489
                           );
   CALCULATION_reg : FD1 port map( D => n6709, CP => CLK_I, Q => n_1037, QN => 
                           n1907);
   v_CALCULATION_CNTR_reg_1_inst : FD1 port map( D => n6652, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_1_port, QN => n367);
   v_CALCULATION_CNTR_reg_2_inst : FD1 port map( D => n6653, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_2_port, QN => n365);
   v_CALCULATION_CNTR_reg_3_inst : FD1 port map( D => n6654, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_3_port, QN => n375);
   v_CALCULATION_CNTR_reg_4_inst : FD1 port map( D => n6655, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_4_port, QN => n317);
   v_CALCULATION_CNTR_reg_5_inst : FD1 port map( D => n8217, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_5_port, QN => n2009);
   v_CALCULATION_CNTR_reg_6_inst : FD1 port map( D => n8218, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_6_port, QN => n2125);
   v_CALCULATION_CNTR_reg_7_inst : FD1 port map( D => n8219, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_7_port, QN => n2006);
   i_INTERN_ADDR_RD0_reg_0_inst : FD1 port map( D => n6708, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD0_0_port, QN => n6649);
   i_INTERN_ADDR_RD0_reg_1_inst : FD1 port map( D => n6707, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD0_1_port, QN => n6648);
   i_INTERN_ADDR_RD0_reg_2_inst : FD1 port map( D => n6706, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD0_2_port, QN => n6647);
   i_INTERN_ADDR_RD0_reg_3_inst : FD1 port map( D => n6705, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD0_3_port, QN => n6646);
   i_INTERN_ADDR_RD0_reg_4_inst : FD1 port map( D => n6704, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD0_4_port, QN => n6645);
   i_INTERN_ADDR_RD0_reg_5_inst : FD1 port map( D => n6703, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD0_5_port, QN => n6644);
   SRAM_WREN0_reg : FD1 port map( D => n6702, CP => CLK_I, Q => n_1038, QN => 
                           n2491);
   i_SRAM_ADDR_WR0_reg_5_inst : FD1 port map( D => n6701, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR0_5_port, QN => n6638);
   i_SRAM_ADDR_WR0_reg_0_inst : FD1 port map( D => n6700, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR0_0_port, QN => n6643);
   i_SRAM_ADDR_WR0_reg_1_inst : FD1 port map( D => n6699, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR0_1_port, QN => n6642);
   i_SRAM_ADDR_WR0_reg_2_inst : FD1 port map( D => n6698, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR0_2_port, QN => n6641);
   i_SRAM_ADDR_WR0_reg_3_inst : FD1 port map( D => n6697, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR0_3_port, QN => n6640);
   i_SRAM_ADDR_WR0_reg_4_inst : FD1 port map( D => n6696, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR0_4_port, QN => n6639);
   v_TEMP_VECTOR_reg_7_inst : FD1 port map( D => n6688, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_7_port, QN => n_1039);
   KEY_EXPAN0_reg_63_7_inst : FD1 port map( D => n5101, CP => CLK_I, Q => 
                           n_1040, QN => n4503);
   KEY_EXPAN0_reg_62_7_inst : FD1 port map( D => n5100, CP => CLK_I, Q => 
                           n_1041, QN => n4502);
   KEY_EXPAN0_reg_61_7_inst : FD1 port map( D => n5099, CP => CLK_I, Q => 
                           n_1042, QN => n4505);
   KEY_EXPAN0_reg_60_7_inst : FD1 port map( D => n5098, CP => CLK_I, Q => 
                           n_1043, QN => n4504);
   KEY_EXPAN0_reg_59_7_inst : FD1 port map( D => n5097, CP => CLK_I, Q => 
                           n_1044, QN => n4507);
   KEY_EXPAN0_reg_58_7_inst : FD1 port map( D => n5096, CP => CLK_I, Q => 
                           n_1045, QN => n4506);
   KEY_EXPAN0_reg_57_7_inst : FD1 port map( D => n5095, CP => CLK_I, Q => 
                           n_1046, QN => n4509);
   KEY_EXPAN0_reg_56_7_inst : FD1 port map( D => n5094, CP => CLK_I, Q => 
                           n_1047, QN => n4508);
   KEY_EXPAN0_reg_55_7_inst : FD1 port map( D => n5093, CP => CLK_I, Q => 
                           n_1048, QN => n4495);
   KEY_EXPAN0_reg_54_7_inst : FD1 port map( D => n5092, CP => CLK_I, Q => 
                           n_1049, QN => n4494);
   KEY_EXPAN0_reg_53_7_inst : FD1 port map( D => n5091, CP => CLK_I, Q => 
                           n_1050, QN => n4497);
   KEY_EXPAN0_reg_52_7_inst : FD1 port map( D => n5090, CP => CLK_I, Q => 
                           n_1051, QN => n4496);
   KEY_EXPAN0_reg_51_7_inst : FD1 port map( D => n5089, CP => CLK_I, Q => 
                           n_1052, QN => n4499);
   KEY_EXPAN0_reg_50_7_inst : FD1 port map( D => n5088, CP => CLK_I, Q => 
                           n_1053, QN => n4498);
   KEY_EXPAN0_reg_49_7_inst : FD1 port map( D => n5087, CP => CLK_I, Q => 
                           n_1054, QN => n4501);
   KEY_EXPAN0_reg_48_7_inst : FD1 port map( D => n5086, CP => CLK_I, Q => 
                           n_1055, QN => n4500);
   KEY_EXPAN0_reg_47_7_inst : FD1 port map( D => n5085, CP => CLK_I, Q => 
                           n_1056, QN => n4487);
   KEY_EXPAN0_reg_46_7_inst : FD1 port map( D => n5084, CP => CLK_I, Q => 
                           n_1057, QN => n4486);
   KEY_EXPAN0_reg_45_7_inst : FD1 port map( D => n5083, CP => CLK_I, Q => 
                           n_1058, QN => n4489);
   KEY_EXPAN0_reg_44_7_inst : FD1 port map( D => n5082, CP => CLK_I, Q => 
                           n_1059, QN => n4488);
   KEY_EXPAN0_reg_43_7_inst : FD1 port map( D => n5081, CP => CLK_I, Q => 
                           n_1060, QN => n4491);
   KEY_EXPAN0_reg_42_7_inst : FD1 port map( D => n5080, CP => CLK_I, Q => 
                           n_1061, QN => n4490);
   KEY_EXPAN0_reg_41_7_inst : FD1 port map( D => n5079, CP => CLK_I, Q => 
                           n_1062, QN => n4493);
   KEY_EXPAN0_reg_40_7_inst : FD1 port map( D => n5078, CP => CLK_I, Q => 
                           n_1063, QN => n4492);
   KEY_EXPAN0_reg_39_7_inst : FD1 port map( D => n5077, CP => CLK_I, Q => 
                           n_1064, QN => n4479);
   KEY_EXPAN0_reg_38_7_inst : FD1 port map( D => n5076, CP => CLK_I, Q => 
                           n_1065, QN => n4478);
   KEY_EXPAN0_reg_37_7_inst : FD1 port map( D => n5075, CP => CLK_I, Q => 
                           n_1066, QN => n4481);
   KEY_EXPAN0_reg_36_7_inst : FD1 port map( D => n5074, CP => CLK_I, Q => 
                           n_1067, QN => n4480);
   KEY_EXPAN0_reg_35_7_inst : FD1 port map( D => n5073, CP => CLK_I, Q => 
                           n_1068, QN => n4483);
   KEY_EXPAN0_reg_34_7_inst : FD1 port map( D => n5072, CP => CLK_I, Q => 
                           n_1069, QN => n4482);
   KEY_EXPAN0_reg_33_7_inst : FD1 port map( D => n5071, CP => CLK_I, Q => 
                           n_1070, QN => n4485);
   KEY_EXPAN0_reg_32_7_inst : FD1 port map( D => n5070, CP => CLK_I, Q => 
                           n_1071, QN => n4484);
   KEY_EXPAN0_reg_31_7_inst : FD1 port map( D => n5069, CP => CLK_I, Q => 
                           n_1072, QN => n4535);
   KEY_EXPAN0_reg_30_7_inst : FD1 port map( D => n5068, CP => CLK_I, Q => 
                           n_1073, QN => n4534);
   KEY_EXPAN0_reg_29_7_inst : FD1 port map( D => n5067, CP => CLK_I, Q => 
                           n_1074, QN => n4537);
   KEY_EXPAN0_reg_28_7_inst : FD1 port map( D => n5066, CP => CLK_I, Q => 
                           n_1075, QN => n4536);
   KEY_EXPAN0_reg_27_7_inst : FD1 port map( D => n5065, CP => CLK_I, Q => 
                           n_1076, QN => n4539);
   KEY_EXPAN0_reg_26_7_inst : FD1 port map( D => n5064, CP => CLK_I, Q => 
                           n_1077, QN => n4538);
   KEY_EXPAN0_reg_25_7_inst : FD1 port map( D => n5063, CP => CLK_I, Q => 
                           n_1078, QN => n4541);
   KEY_EXPAN0_reg_24_7_inst : FD1 port map( D => n5062, CP => CLK_I, Q => 
                           n_1079, QN => n4540);
   KEY_EXPAN0_reg_23_7_inst : FD1 port map( D => n5061, CP => CLK_I, Q => 
                           n_1080, QN => n4527);
   KEY_EXPAN0_reg_22_7_inst : FD1 port map( D => n5060, CP => CLK_I, Q => 
                           n_1081, QN => n4526);
   KEY_EXPAN0_reg_21_7_inst : FD1 port map( D => n5059, CP => CLK_I, Q => 
                           n_1082, QN => n4529);
   KEY_EXPAN0_reg_20_7_inst : FD1 port map( D => n5058, CP => CLK_I, Q => 
                           n_1083, QN => n4528);
   KEY_EXPAN0_reg_19_7_inst : FD1 port map( D => n5057, CP => CLK_I, Q => 
                           n_1084, QN => n4531);
   KEY_EXPAN0_reg_18_7_inst : FD1 port map( D => n5056, CP => CLK_I, Q => 
                           n_1085, QN => n4530);
   KEY_EXPAN0_reg_17_7_inst : FD1 port map( D => n5055, CP => CLK_I, Q => 
                           n_1086, QN => n4533);
   KEY_EXPAN0_reg_16_7_inst : FD1 port map( D => n5054, CP => CLK_I, Q => 
                           n_1087, QN => n4532);
   KEY_EXPAN0_reg_15_7_inst : FD1 port map( D => n5053, CP => CLK_I, Q => 
                           n_1088, QN => n4519);
   KEY_EXPAN0_reg_14_7_inst : FD1 port map( D => n5052, CP => CLK_I, Q => 
                           n_1089, QN => n4518);
   KEY_EXPAN0_reg_13_7_inst : FD1 port map( D => n5051, CP => CLK_I, Q => 
                           n_1090, QN => n4521);
   KEY_EXPAN0_reg_12_7_inst : FD1 port map( D => n5050, CP => CLK_I, Q => 
                           n_1091, QN => n4520);
   KEY_EXPAN0_reg_11_7_inst : FD1 port map( D => n5049, CP => CLK_I, Q => 
                           n_1092, QN => n4523);
   KEY_EXPAN0_reg_10_7_inst : FD1 port map( D => n5048, CP => CLK_I, Q => 
                           n_1093, QN => n4522);
   KEY_EXPAN0_reg_9_7_inst : FD1 port map( D => n5047, CP => CLK_I, Q => n_1094
                           , QN => n4525);
   KEY_EXPAN0_reg_8_7_inst : FD1 port map( D => n5046, CP => CLK_I, Q => n_1095
                           , QN => n4524);
   KEY_EXPAN0_reg_7_7_inst : FD1 port map( D => n5045, CP => CLK_I, Q => n_1096
                           , QN => n4511);
   KEY_EXPAN0_reg_6_7_inst : FD1 port map( D => n5044, CP => CLK_I, Q => n_1097
                           , QN => n4510);
   KEY_EXPAN0_reg_5_7_inst : FD1 port map( D => n5043, CP => CLK_I, Q => n_1098
                           , QN => n4513);
   KEY_EXPAN0_reg_4_7_inst : FD1 port map( D => n5042, CP => CLK_I, Q => n_1099
                           , QN => n4512);
   KEY_EXPAN0_reg_3_7_inst : FD1 port map( D => n5041, CP => CLK_I, Q => n_1100
                           , QN => n4515);
   KEY_EXPAN0_reg_2_7_inst : FD1 port map( D => n5040, CP => CLK_I, Q => n_1101
                           , QN => n4514);
   KEY_EXPAN0_reg_1_7_inst : FD1 port map( D => n5039, CP => CLK_I, Q => n_1102
                           , QN => n4517);
   KEY_EXPAN0_reg_0_7_inst : FD1 port map( D => n5038, CP => CLK_I, Q => n_1103
                           , QN => n4516);
   v_KEY_COL_OUT0_reg_7_inst : FD1 port map( D => n4580, CP => CLK_I, Q => 
                           n_1104, QN => n354);
   v_TEMP_VECTOR_reg_31_inst : FD1 port map( D => n6664, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_31_port, QN => n_1105);
   KEY_EXPAN0_reg_63_31_inst : FD1 port map( D => n6637, CP => CLK_I, Q => 
                           n_1106, QN => n4439);
   KEY_EXPAN0_reg_62_31_inst : FD1 port map( D => n6636, CP => CLK_I, Q => 
                           n_1107, QN => n4438);
   KEY_EXPAN0_reg_61_31_inst : FD1 port map( D => n6635, CP => CLK_I, Q => 
                           n_1108, QN => n4441);
   KEY_EXPAN0_reg_60_31_inst : FD1 port map( D => n6634, CP => CLK_I, Q => 
                           n_1109, QN => n4440);
   KEY_EXPAN0_reg_59_31_inst : FD1 port map( D => n6633, CP => CLK_I, Q => 
                           n_1110, QN => n4443);
   KEY_EXPAN0_reg_58_31_inst : FD1 port map( D => n6632, CP => CLK_I, Q => 
                           n_1111, QN => n4442);
   KEY_EXPAN0_reg_57_31_inst : FD1 port map( D => n6631, CP => CLK_I, Q => 
                           n_1112, QN => n4445);
   KEY_EXPAN0_reg_56_31_inst : FD1 port map( D => n6630, CP => CLK_I, Q => 
                           n_1113, QN => n4444);
   KEY_EXPAN0_reg_55_31_inst : FD1 port map( D => n6629, CP => CLK_I, Q => 
                           n_1114, QN => n4431);
   KEY_EXPAN0_reg_54_31_inst : FD1 port map( D => n6628, CP => CLK_I, Q => 
                           n_1115, QN => n4430);
   KEY_EXPAN0_reg_53_31_inst : FD1 port map( D => n6627, CP => CLK_I, Q => 
                           n_1116, QN => n4433);
   KEY_EXPAN0_reg_52_31_inst : FD1 port map( D => n6626, CP => CLK_I, Q => 
                           n_1117, QN => n4432);
   KEY_EXPAN0_reg_51_31_inst : FD1 port map( D => n6625, CP => CLK_I, Q => 
                           n_1118, QN => n4435);
   KEY_EXPAN0_reg_50_31_inst : FD1 port map( D => n6624, CP => CLK_I, Q => 
                           n_1119, QN => n4434);
   KEY_EXPAN0_reg_49_31_inst : FD1 port map( D => n6623, CP => CLK_I, Q => 
                           n_1120, QN => n4437);
   KEY_EXPAN0_reg_48_31_inst : FD1 port map( D => n6622, CP => CLK_I, Q => 
                           n_1121, QN => n4436);
   KEY_EXPAN0_reg_47_31_inst : FD1 port map( D => n6621, CP => CLK_I, Q => 
                           n_1122, QN => n4423);
   KEY_EXPAN0_reg_46_31_inst : FD1 port map( D => n6620, CP => CLK_I, Q => 
                           n_1123, QN => n4422);
   KEY_EXPAN0_reg_45_31_inst : FD1 port map( D => n6619, CP => CLK_I, Q => 
                           n_1124, QN => n4425);
   KEY_EXPAN0_reg_44_31_inst : FD1 port map( D => n6618, CP => CLK_I, Q => 
                           n_1125, QN => n4424);
   KEY_EXPAN0_reg_43_31_inst : FD1 port map( D => n6617, CP => CLK_I, Q => 
                           n_1126, QN => n4427);
   KEY_EXPAN0_reg_42_31_inst : FD1 port map( D => n6616, CP => CLK_I, Q => 
                           n_1127, QN => n4426);
   KEY_EXPAN0_reg_41_31_inst : FD1 port map( D => n6615, CP => CLK_I, Q => 
                           n_1128, QN => n4429);
   KEY_EXPAN0_reg_40_31_inst : FD1 port map( D => n6614, CP => CLK_I, Q => 
                           n_1129, QN => n4428);
   KEY_EXPAN0_reg_39_31_inst : FD1 port map( D => n6613, CP => CLK_I, Q => 
                           n_1130, QN => n4415);
   KEY_EXPAN0_reg_38_31_inst : FD1 port map( D => n6612, CP => CLK_I, Q => 
                           n_1131, QN => n4414);
   KEY_EXPAN0_reg_37_31_inst : FD1 port map( D => n6611, CP => CLK_I, Q => 
                           n_1132, QN => n4417);
   KEY_EXPAN0_reg_36_31_inst : FD1 port map( D => n6610, CP => CLK_I, Q => 
                           n_1133, QN => n4416);
   KEY_EXPAN0_reg_35_31_inst : FD1 port map( D => n6609, CP => CLK_I, Q => 
                           n_1134, QN => n4419);
   KEY_EXPAN0_reg_34_31_inst : FD1 port map( D => n6608, CP => CLK_I, Q => 
                           n_1135, QN => n4418);
   KEY_EXPAN0_reg_33_31_inst : FD1 port map( D => n6607, CP => CLK_I, Q => 
                           n_1136, QN => n4421);
   KEY_EXPAN0_reg_32_31_inst : FD1 port map( D => n6606, CP => CLK_I, Q => 
                           n_1137, QN => n4420);
   KEY_EXPAN0_reg_31_31_inst : FD1 port map( D => n6605, CP => CLK_I, Q => 
                           n_1138, QN => n4471);
   KEY_EXPAN0_reg_30_31_inst : FD1 port map( D => n6604, CP => CLK_I, Q => 
                           n_1139, QN => n4470);
   KEY_EXPAN0_reg_29_31_inst : FD1 port map( D => n6603, CP => CLK_I, Q => 
                           n_1140, QN => n4473);
   KEY_EXPAN0_reg_28_31_inst : FD1 port map( D => n6602, CP => CLK_I, Q => 
                           n_1141, QN => n4472);
   KEY_EXPAN0_reg_27_31_inst : FD1 port map( D => n6601, CP => CLK_I, Q => 
                           n_1142, QN => n4475);
   KEY_EXPAN0_reg_26_31_inst : FD1 port map( D => n6600, CP => CLK_I, Q => 
                           n_1143, QN => n4474);
   KEY_EXPAN0_reg_25_31_inst : FD1 port map( D => n6599, CP => CLK_I, Q => 
                           n_1144, QN => n4477);
   KEY_EXPAN0_reg_24_31_inst : FD1 port map( D => n6598, CP => CLK_I, Q => 
                           n_1145, QN => n4476);
   KEY_EXPAN0_reg_23_31_inst : FD1 port map( D => n6597, CP => CLK_I, Q => 
                           n_1146, QN => n4463);
   KEY_EXPAN0_reg_22_31_inst : FD1 port map( D => n6596, CP => CLK_I, Q => 
                           n_1147, QN => n4462);
   KEY_EXPAN0_reg_21_31_inst : FD1 port map( D => n6595, CP => CLK_I, Q => 
                           n_1148, QN => n4465);
   KEY_EXPAN0_reg_20_31_inst : FD1 port map( D => n6594, CP => CLK_I, Q => 
                           n_1149, QN => n4464);
   KEY_EXPAN0_reg_19_31_inst : FD1 port map( D => n6593, CP => CLK_I, Q => 
                           n_1150, QN => n4467);
   KEY_EXPAN0_reg_18_31_inst : FD1 port map( D => n6592, CP => CLK_I, Q => 
                           n_1151, QN => n4466);
   KEY_EXPAN0_reg_17_31_inst : FD1 port map( D => n6591, CP => CLK_I, Q => 
                           n_1152, QN => n4469);
   KEY_EXPAN0_reg_16_31_inst : FD1 port map( D => n6590, CP => CLK_I, Q => 
                           n_1153, QN => n4468);
   KEY_EXPAN0_reg_15_31_inst : FD1 port map( D => n6589, CP => CLK_I, Q => 
                           n_1154, QN => n4455);
   KEY_EXPAN0_reg_14_31_inst : FD1 port map( D => n6588, CP => CLK_I, Q => 
                           n_1155, QN => n4454);
   KEY_EXPAN0_reg_13_31_inst : FD1 port map( D => n6587, CP => CLK_I, Q => 
                           n_1156, QN => n4457);
   KEY_EXPAN0_reg_12_31_inst : FD1 port map( D => n6586, CP => CLK_I, Q => 
                           n_1157, QN => n4456);
   KEY_EXPAN0_reg_11_31_inst : FD1 port map( D => n6585, CP => CLK_I, Q => 
                           n_1158, QN => n4459);
   KEY_EXPAN0_reg_10_31_inst : FD1 port map( D => n6584, CP => CLK_I, Q => 
                           n_1159, QN => n4458);
   KEY_EXPAN0_reg_9_31_inst : FD1 port map( D => n6583, CP => CLK_I, Q => 
                           n_1160, QN => n4461);
   KEY_EXPAN0_reg_8_31_inst : FD1 port map( D => n6582, CP => CLK_I, Q => 
                           n_1161, QN => n4460);
   KEY_EXPAN0_reg_7_31_inst : FD1 port map( D => n6581, CP => CLK_I, Q => 
                           n_1162, QN => n4447);
   KEY_EXPAN0_reg_6_31_inst : FD1 port map( D => n6580, CP => CLK_I, Q => 
                           n_1163, QN => n4446);
   KEY_EXPAN0_reg_5_31_inst : FD1 port map( D => n6579, CP => CLK_I, Q => 
                           n_1164, QN => n4449);
   KEY_EXPAN0_reg_4_31_inst : FD1 port map( D => n6578, CP => CLK_I, Q => 
                           n_1165, QN => n4448);
   KEY_EXPAN0_reg_3_31_inst : FD1 port map( D => n6577, CP => CLK_I, Q => 
                           n_1166, QN => n4451);
   KEY_EXPAN0_reg_2_31_inst : FD1 port map( D => n6576, CP => CLK_I, Q => 
                           n_1167, QN => n4450);
   KEY_EXPAN0_reg_1_31_inst : FD1 port map( D => n6575, CP => CLK_I, Q => 
                           n_1168, QN => n4453);
   KEY_EXPAN0_reg_0_31_inst : FD1 port map( D => n6574, CP => CLK_I, Q => 
                           n_1169, QN => n4452);
   v_KEY_COL_OUT0_reg_31_inst : FD1 port map( D => n4579, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_31_port, QN => n1498);
   v_TEMP_VECTOR_reg_23_inst : FD1 port map( D => n6672, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_23_port, QN => n_1170);
   KEY_EXPAN0_reg_63_23_inst : FD1 port map( D => n6125, CP => CLK_I, Q => 
                           n_1171, QN => n4375);
   KEY_EXPAN0_reg_62_23_inst : FD1 port map( D => n6124, CP => CLK_I, Q => 
                           n_1172, QN => n4374);
   KEY_EXPAN0_reg_61_23_inst : FD1 port map( D => n6123, CP => CLK_I, Q => 
                           n_1173, QN => n4377);
   KEY_EXPAN0_reg_60_23_inst : FD1 port map( D => n6122, CP => CLK_I, Q => 
                           n_1174, QN => n4376);
   KEY_EXPAN0_reg_59_23_inst : FD1 port map( D => n6121, CP => CLK_I, Q => 
                           n_1175, QN => n4379);
   KEY_EXPAN0_reg_58_23_inst : FD1 port map( D => n6120, CP => CLK_I, Q => 
                           n_1176, QN => n4378);
   KEY_EXPAN0_reg_57_23_inst : FD1 port map( D => n6119, CP => CLK_I, Q => 
                           n_1177, QN => n4381);
   KEY_EXPAN0_reg_56_23_inst : FD1 port map( D => n6118, CP => CLK_I, Q => 
                           n_1178, QN => n4380);
   KEY_EXPAN0_reg_55_23_inst : FD1 port map( D => n6117, CP => CLK_I, Q => 
                           n_1179, QN => n4367);
   KEY_EXPAN0_reg_54_23_inst : FD1 port map( D => n6116, CP => CLK_I, Q => 
                           n_1180, QN => n4366);
   KEY_EXPAN0_reg_53_23_inst : FD1 port map( D => n6115, CP => CLK_I, Q => 
                           n_1181, QN => n4369);
   KEY_EXPAN0_reg_52_23_inst : FD1 port map( D => n6114, CP => CLK_I, Q => 
                           n_1182, QN => n4368);
   KEY_EXPAN0_reg_51_23_inst : FD1 port map( D => n6113, CP => CLK_I, Q => 
                           n_1183, QN => n4371);
   KEY_EXPAN0_reg_50_23_inst : FD1 port map( D => n6112, CP => CLK_I, Q => 
                           n_1184, QN => n4370);
   KEY_EXPAN0_reg_49_23_inst : FD1 port map( D => n6111, CP => CLK_I, Q => 
                           n_1185, QN => n4373);
   KEY_EXPAN0_reg_48_23_inst : FD1 port map( D => n6110, CP => CLK_I, Q => 
                           n_1186, QN => n4372);
   KEY_EXPAN0_reg_47_23_inst : FD1 port map( D => n6109, CP => CLK_I, Q => 
                           n_1187, QN => n4359);
   KEY_EXPAN0_reg_46_23_inst : FD1 port map( D => n6108, CP => CLK_I, Q => 
                           n_1188, QN => n4358);
   KEY_EXPAN0_reg_45_23_inst : FD1 port map( D => n6107, CP => CLK_I, Q => 
                           n_1189, QN => n4361);
   KEY_EXPAN0_reg_44_23_inst : FD1 port map( D => n6106, CP => CLK_I, Q => 
                           n_1190, QN => n4360);
   KEY_EXPAN0_reg_43_23_inst : FD1 port map( D => n6105, CP => CLK_I, Q => 
                           n_1191, QN => n4363);
   KEY_EXPAN0_reg_42_23_inst : FD1 port map( D => n6104, CP => CLK_I, Q => 
                           n_1192, QN => n4362);
   KEY_EXPAN0_reg_41_23_inst : FD1 port map( D => n6103, CP => CLK_I, Q => 
                           n_1193, QN => n4365);
   KEY_EXPAN0_reg_40_23_inst : FD1 port map( D => n6102, CP => CLK_I, Q => 
                           n_1194, QN => n4364);
   KEY_EXPAN0_reg_39_23_inst : FD1 port map( D => n6101, CP => CLK_I, Q => 
                           n_1195, QN => n4351);
   KEY_EXPAN0_reg_38_23_inst : FD1 port map( D => n6100, CP => CLK_I, Q => 
                           n_1196, QN => n4350);
   KEY_EXPAN0_reg_37_23_inst : FD1 port map( D => n6099, CP => CLK_I, Q => 
                           n_1197, QN => n4353);
   KEY_EXPAN0_reg_36_23_inst : FD1 port map( D => n6098, CP => CLK_I, Q => 
                           n_1198, QN => n4352);
   KEY_EXPAN0_reg_35_23_inst : FD1 port map( D => n6097, CP => CLK_I, Q => 
                           n_1199, QN => n4355);
   KEY_EXPAN0_reg_34_23_inst : FD1 port map( D => n6096, CP => CLK_I, Q => 
                           n_1200, QN => n4354);
   KEY_EXPAN0_reg_33_23_inst : FD1 port map( D => n6095, CP => CLK_I, Q => 
                           n_1201, QN => n4357);
   KEY_EXPAN0_reg_32_23_inst : FD1 port map( D => n6094, CP => CLK_I, Q => 
                           n_1202, QN => n4356);
   KEY_EXPAN0_reg_31_23_inst : FD1 port map( D => n6093, CP => CLK_I, Q => 
                           n_1203, QN => n4407);
   KEY_EXPAN0_reg_30_23_inst : FD1 port map( D => n6092, CP => CLK_I, Q => 
                           n_1204, QN => n4406);
   KEY_EXPAN0_reg_29_23_inst : FD1 port map( D => n6091, CP => CLK_I, Q => 
                           n_1205, QN => n4409);
   KEY_EXPAN0_reg_28_23_inst : FD1 port map( D => n6090, CP => CLK_I, Q => 
                           n_1206, QN => n4408);
   KEY_EXPAN0_reg_27_23_inst : FD1 port map( D => n6089, CP => CLK_I, Q => 
                           n_1207, QN => n4411);
   KEY_EXPAN0_reg_26_23_inst : FD1 port map( D => n6088, CP => CLK_I, Q => 
                           n_1208, QN => n4410);
   KEY_EXPAN0_reg_25_23_inst : FD1 port map( D => n6087, CP => CLK_I, Q => 
                           n_1209, QN => n4413);
   KEY_EXPAN0_reg_24_23_inst : FD1 port map( D => n6086, CP => CLK_I, Q => 
                           n_1210, QN => n4412);
   KEY_EXPAN0_reg_23_23_inst : FD1 port map( D => n6085, CP => CLK_I, Q => 
                           n_1211, QN => n4399);
   KEY_EXPAN0_reg_22_23_inst : FD1 port map( D => n6084, CP => CLK_I, Q => 
                           n_1212, QN => n4398);
   KEY_EXPAN0_reg_21_23_inst : FD1 port map( D => n6083, CP => CLK_I, Q => 
                           n_1213, QN => n4401);
   KEY_EXPAN0_reg_20_23_inst : FD1 port map( D => n6082, CP => CLK_I, Q => 
                           n_1214, QN => n4400);
   KEY_EXPAN0_reg_19_23_inst : FD1 port map( D => n6081, CP => CLK_I, Q => 
                           n_1215, QN => n4403);
   KEY_EXPAN0_reg_18_23_inst : FD1 port map( D => n6080, CP => CLK_I, Q => 
                           n_1216, QN => n4402);
   KEY_EXPAN0_reg_17_23_inst : FD1 port map( D => n6079, CP => CLK_I, Q => 
                           n_1217, QN => n4405);
   KEY_EXPAN0_reg_16_23_inst : FD1 port map( D => n6078, CP => CLK_I, Q => 
                           n_1218, QN => n4404);
   KEY_EXPAN0_reg_15_23_inst : FD1 port map( D => n6077, CP => CLK_I, Q => 
                           n_1219, QN => n4391);
   KEY_EXPAN0_reg_14_23_inst : FD1 port map( D => n6076, CP => CLK_I, Q => 
                           n_1220, QN => n4390);
   KEY_EXPAN0_reg_13_23_inst : FD1 port map( D => n6075, CP => CLK_I, Q => 
                           n_1221, QN => n4393);
   KEY_EXPAN0_reg_12_23_inst : FD1 port map( D => n6074, CP => CLK_I, Q => 
                           n_1222, QN => n4392);
   KEY_EXPAN0_reg_11_23_inst : FD1 port map( D => n6073, CP => CLK_I, Q => 
                           n_1223, QN => n4395);
   KEY_EXPAN0_reg_10_23_inst : FD1 port map( D => n6072, CP => CLK_I, Q => 
                           n_1224, QN => n4394);
   KEY_EXPAN0_reg_9_23_inst : FD1 port map( D => n6071, CP => CLK_I, Q => 
                           n_1225, QN => n4397);
   KEY_EXPAN0_reg_8_23_inst : FD1 port map( D => n6070, CP => CLK_I, Q => 
                           n_1226, QN => n4396);
   KEY_EXPAN0_reg_7_23_inst : FD1 port map( D => n6069, CP => CLK_I, Q => 
                           n_1227, QN => n4383);
   KEY_EXPAN0_reg_6_23_inst : FD1 port map( D => n6068, CP => CLK_I, Q => 
                           n_1228, QN => n4382);
   KEY_EXPAN0_reg_5_23_inst : FD1 port map( D => n6067, CP => CLK_I, Q => 
                           n_1229, QN => n4385);
   KEY_EXPAN0_reg_4_23_inst : FD1 port map( D => n6066, CP => CLK_I, Q => 
                           n_1230, QN => n4384);
   KEY_EXPAN0_reg_3_23_inst : FD1 port map( D => n6065, CP => CLK_I, Q => 
                           n_1231, QN => n4387);
   KEY_EXPAN0_reg_2_23_inst : FD1 port map( D => n6064, CP => CLK_I, Q => 
                           n_1232, QN => n4386);
   KEY_EXPAN0_reg_1_23_inst : FD1 port map( D => n6063, CP => CLK_I, Q => 
                           n_1233, QN => n4389);
   KEY_EXPAN0_reg_0_23_inst : FD1 port map( D => n6062, CP => CLK_I, Q => 
                           n_1234, QN => n4388);
   v_KEY_COL_OUT0_reg_23_inst : FD1 port map( D => n4578, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_23_port, QN => n390);
   v_TEMP_VECTOR_reg_15_inst : FD1 port map( D => n6680, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_15_port, QN => n_1235);
   KEY_EXPAN0_reg_63_15_inst : FD1 port map( D => n5613, CP => CLK_I, Q => 
                           n_1236, QN => n4311);
   KEY_EXPAN0_reg_62_15_inst : FD1 port map( D => n5612, CP => CLK_I, Q => 
                           n_1237, QN => n4310);
   KEY_EXPAN0_reg_61_15_inst : FD1 port map( D => n5611, CP => CLK_I, Q => 
                           n_1238, QN => n4313);
   KEY_EXPAN0_reg_60_15_inst : FD1 port map( D => n5610, CP => CLK_I, Q => 
                           n_1239, QN => n4312);
   KEY_EXPAN0_reg_59_15_inst : FD1 port map( D => n5609, CP => CLK_I, Q => 
                           n_1240, QN => n4315);
   KEY_EXPAN0_reg_58_15_inst : FD1 port map( D => n5608, CP => CLK_I, Q => 
                           n_1241, QN => n4314);
   KEY_EXPAN0_reg_57_15_inst : FD1 port map( D => n5607, CP => CLK_I, Q => 
                           n_1242, QN => n4317);
   KEY_EXPAN0_reg_56_15_inst : FD1 port map( D => n5606, CP => CLK_I, Q => 
                           n_1243, QN => n4316);
   KEY_EXPAN0_reg_55_15_inst : FD1 port map( D => n5605, CP => CLK_I, Q => 
                           n_1244, QN => n4303);
   KEY_EXPAN0_reg_54_15_inst : FD1 port map( D => n5604, CP => CLK_I, Q => 
                           n_1245, QN => n4302);
   KEY_EXPAN0_reg_53_15_inst : FD1 port map( D => n5603, CP => CLK_I, Q => 
                           n_1246, QN => n4305);
   KEY_EXPAN0_reg_52_15_inst : FD1 port map( D => n5602, CP => CLK_I, Q => 
                           n_1247, QN => n4304);
   KEY_EXPAN0_reg_51_15_inst : FD1 port map( D => n5601, CP => CLK_I, Q => 
                           n_1248, QN => n4307);
   KEY_EXPAN0_reg_50_15_inst : FD1 port map( D => n5600, CP => CLK_I, Q => 
                           n_1249, QN => n4306);
   KEY_EXPAN0_reg_49_15_inst : FD1 port map( D => n5599, CP => CLK_I, Q => 
                           n_1250, QN => n4309);
   KEY_EXPAN0_reg_48_15_inst : FD1 port map( D => n5598, CP => CLK_I, Q => 
                           n_1251, QN => n4308);
   KEY_EXPAN0_reg_47_15_inst : FD1 port map( D => n5597, CP => CLK_I, Q => 
                           n_1252, QN => n4295);
   KEY_EXPAN0_reg_46_15_inst : FD1 port map( D => n5596, CP => CLK_I, Q => 
                           n_1253, QN => n4294);
   KEY_EXPAN0_reg_45_15_inst : FD1 port map( D => n5595, CP => CLK_I, Q => 
                           n_1254, QN => n4297);
   KEY_EXPAN0_reg_44_15_inst : FD1 port map( D => n5594, CP => CLK_I, Q => 
                           n_1255, QN => n4296);
   KEY_EXPAN0_reg_43_15_inst : FD1 port map( D => n5593, CP => CLK_I, Q => 
                           n_1256, QN => n4299);
   KEY_EXPAN0_reg_42_15_inst : FD1 port map( D => n5592, CP => CLK_I, Q => 
                           n_1257, QN => n4298);
   KEY_EXPAN0_reg_41_15_inst : FD1 port map( D => n5591, CP => CLK_I, Q => 
                           n_1258, QN => n4301);
   KEY_EXPAN0_reg_40_15_inst : FD1 port map( D => n5590, CP => CLK_I, Q => 
                           n_1259, QN => n4300);
   KEY_EXPAN0_reg_39_15_inst : FD1 port map( D => n5589, CP => CLK_I, Q => 
                           n_1260, QN => n4287);
   KEY_EXPAN0_reg_38_15_inst : FD1 port map( D => n5588, CP => CLK_I, Q => 
                           n_1261, QN => n4286);
   KEY_EXPAN0_reg_37_15_inst : FD1 port map( D => n5587, CP => CLK_I, Q => 
                           n_1262, QN => n4289);
   KEY_EXPAN0_reg_36_15_inst : FD1 port map( D => n5586, CP => CLK_I, Q => 
                           n_1263, QN => n4288);
   KEY_EXPAN0_reg_35_15_inst : FD1 port map( D => n5585, CP => CLK_I, Q => 
                           n_1264, QN => n4291);
   KEY_EXPAN0_reg_34_15_inst : FD1 port map( D => n5584, CP => CLK_I, Q => 
                           n_1265, QN => n4290);
   KEY_EXPAN0_reg_33_15_inst : FD1 port map( D => n5583, CP => CLK_I, Q => 
                           n_1266, QN => n4293);
   KEY_EXPAN0_reg_32_15_inst : FD1 port map( D => n5582, CP => CLK_I, Q => 
                           n_1267, QN => n4292);
   KEY_EXPAN0_reg_31_15_inst : FD1 port map( D => n5581, CP => CLK_I, Q => 
                           n_1268, QN => n4343);
   KEY_EXPAN0_reg_30_15_inst : FD1 port map( D => n5580, CP => CLK_I, Q => 
                           n_1269, QN => n4342);
   KEY_EXPAN0_reg_29_15_inst : FD1 port map( D => n5579, CP => CLK_I, Q => 
                           n_1270, QN => n4345);
   KEY_EXPAN0_reg_28_15_inst : FD1 port map( D => n5578, CP => CLK_I, Q => 
                           n_1271, QN => n4344);
   KEY_EXPAN0_reg_27_15_inst : FD1 port map( D => n5577, CP => CLK_I, Q => 
                           n_1272, QN => n4347);
   KEY_EXPAN0_reg_26_15_inst : FD1 port map( D => n5576, CP => CLK_I, Q => 
                           n_1273, QN => n4346);
   KEY_EXPAN0_reg_25_15_inst : FD1 port map( D => n5575, CP => CLK_I, Q => 
                           n_1274, QN => n4349);
   KEY_EXPAN0_reg_24_15_inst : FD1 port map( D => n5574, CP => CLK_I, Q => 
                           n_1275, QN => n4348);
   KEY_EXPAN0_reg_23_15_inst : FD1 port map( D => n5573, CP => CLK_I, Q => 
                           n_1276, QN => n4335);
   KEY_EXPAN0_reg_22_15_inst : FD1 port map( D => n5572, CP => CLK_I, Q => 
                           n_1277, QN => n4334);
   KEY_EXPAN0_reg_21_15_inst : FD1 port map( D => n5571, CP => CLK_I, Q => 
                           n_1278, QN => n4337);
   KEY_EXPAN0_reg_20_15_inst : FD1 port map( D => n5570, CP => CLK_I, Q => 
                           n_1279, QN => n4336);
   KEY_EXPAN0_reg_19_15_inst : FD1 port map( D => n5569, CP => CLK_I, Q => 
                           n_1280, QN => n4339);
   KEY_EXPAN0_reg_18_15_inst : FD1 port map( D => n5568, CP => CLK_I, Q => 
                           n_1281, QN => n4338);
   KEY_EXPAN0_reg_17_15_inst : FD1 port map( D => n5567, CP => CLK_I, Q => 
                           n_1282, QN => n4341);
   KEY_EXPAN0_reg_16_15_inst : FD1 port map( D => n5566, CP => CLK_I, Q => 
                           n_1283, QN => n4340);
   KEY_EXPAN0_reg_15_15_inst : FD1 port map( D => n5565, CP => CLK_I, Q => 
                           n_1284, QN => n4327);
   KEY_EXPAN0_reg_14_15_inst : FD1 port map( D => n5564, CP => CLK_I, Q => 
                           n_1285, QN => n4326);
   KEY_EXPAN0_reg_13_15_inst : FD1 port map( D => n5563, CP => CLK_I, Q => 
                           n_1286, QN => n4329);
   KEY_EXPAN0_reg_12_15_inst : FD1 port map( D => n5562, CP => CLK_I, Q => 
                           n_1287, QN => n4328);
   KEY_EXPAN0_reg_11_15_inst : FD1 port map( D => n5561, CP => CLK_I, Q => 
                           n_1288, QN => n4331);
   KEY_EXPAN0_reg_10_15_inst : FD1 port map( D => n5560, CP => CLK_I, Q => 
                           n_1289, QN => n4330);
   KEY_EXPAN0_reg_9_15_inst : FD1 port map( D => n5559, CP => CLK_I, Q => 
                           n_1290, QN => n4333);
   KEY_EXPAN0_reg_8_15_inst : FD1 port map( D => n5558, CP => CLK_I, Q => 
                           n_1291, QN => n4332);
   KEY_EXPAN0_reg_7_15_inst : FD1 port map( D => n5557, CP => CLK_I, Q => 
                           n_1292, QN => n4319);
   KEY_EXPAN0_reg_6_15_inst : FD1 port map( D => n5556, CP => CLK_I, Q => 
                           n_1293, QN => n4318);
   KEY_EXPAN0_reg_5_15_inst : FD1 port map( D => n5555, CP => CLK_I, Q => 
                           n_1294, QN => n4321);
   KEY_EXPAN0_reg_4_15_inst : FD1 port map( D => n5554, CP => CLK_I, Q => 
                           n_1295, QN => n4320);
   KEY_EXPAN0_reg_3_15_inst : FD1 port map( D => n5553, CP => CLK_I, Q => 
                           n_1296, QN => n4323);
   KEY_EXPAN0_reg_2_15_inst : FD1 port map( D => n5552, CP => CLK_I, Q => 
                           n_1297, QN => n4322);
   KEY_EXPAN0_reg_1_15_inst : FD1 port map( D => n5551, CP => CLK_I, Q => 
                           n_1298, QN => n4325);
   KEY_EXPAN0_reg_0_15_inst : FD1 port map( D => n5550, CP => CLK_I, Q => 
                           n_1299, QN => n4324);
   v_KEY_COL_OUT0_reg_15_inst : FD1 port map( D => n4577, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_15_port, QN => n387);
   v_TEMP_VECTOR_reg_6_inst : FD1 port map( D => n6689, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_6_port, QN => n2004);
   KEY_EXPAN0_reg_63_6_inst : FD1 port map( D => n5037, CP => CLK_I, Q => 
                           n_1300, QN => n4246);
   KEY_EXPAN0_reg_62_6_inst : FD1 port map( D => n5036, CP => CLK_I, Q => 
                           n_1301, QN => n4245);
   KEY_EXPAN0_reg_61_6_inst : FD1 port map( D => n5035, CP => CLK_I, Q => 
                           n_1302, QN => n4248);
   KEY_EXPAN0_reg_60_6_inst : FD1 port map( D => n5034, CP => CLK_I, Q => 
                           n_1303, QN => n4247);
   KEY_EXPAN0_reg_59_6_inst : FD1 port map( D => n5033, CP => CLK_I, Q => 
                           n_1304, QN => n4250);
   KEY_EXPAN0_reg_58_6_inst : FD1 port map( D => n5032, CP => CLK_I, Q => 
                           n_1305, QN => n4249);
   KEY_EXPAN0_reg_57_6_inst : FD1 port map( D => n5031, CP => CLK_I, Q => 
                           n_1306, QN => n4252);
   KEY_EXPAN0_reg_56_6_inst : FD1 port map( D => n5030, CP => CLK_I, Q => 
                           n_1307, QN => n4251);
   KEY_EXPAN0_reg_55_6_inst : FD1 port map( D => n5029, CP => CLK_I, Q => 
                           n_1308, QN => n4238);
   KEY_EXPAN0_reg_54_6_inst : FD1 port map( D => n5028, CP => CLK_I, Q => 
                           n_1309, QN => n4237);
   KEY_EXPAN0_reg_53_6_inst : FD1 port map( D => n5027, CP => CLK_I, Q => 
                           n_1310, QN => n4240);
   KEY_EXPAN0_reg_52_6_inst : FD1 port map( D => n5026, CP => CLK_I, Q => 
                           n_1311, QN => n4239);
   KEY_EXPAN0_reg_51_6_inst : FD1 port map( D => n5025, CP => CLK_I, Q => 
                           n_1312, QN => n4242);
   KEY_EXPAN0_reg_50_6_inst : FD1 port map( D => n5024, CP => CLK_I, Q => 
                           n_1313, QN => n4241);
   KEY_EXPAN0_reg_49_6_inst : FD1 port map( D => n5023, CP => CLK_I, Q => 
                           n_1314, QN => n4244);
   KEY_EXPAN0_reg_48_6_inst : FD1 port map( D => n5022, CP => CLK_I, Q => 
                           n_1315, QN => n4243);
   KEY_EXPAN0_reg_47_6_inst : FD1 port map( D => n5021, CP => CLK_I, Q => 
                           n_1316, QN => n4230);
   KEY_EXPAN0_reg_46_6_inst : FD1 port map( D => n5020, CP => CLK_I, Q => 
                           n_1317, QN => n4229);
   KEY_EXPAN0_reg_45_6_inst : FD1 port map( D => n5019, CP => CLK_I, Q => 
                           n_1318, QN => n4232);
   KEY_EXPAN0_reg_44_6_inst : FD1 port map( D => n5018, CP => CLK_I, Q => 
                           n_1319, QN => n4231);
   KEY_EXPAN0_reg_43_6_inst : FD1 port map( D => n5017, CP => CLK_I, Q => 
                           n_1320, QN => n4234);
   KEY_EXPAN0_reg_42_6_inst : FD1 port map( D => n5016, CP => CLK_I, Q => 
                           n_1321, QN => n4233);
   KEY_EXPAN0_reg_41_6_inst : FD1 port map( D => n5015, CP => CLK_I, Q => 
                           n_1322, QN => n4236);
   KEY_EXPAN0_reg_40_6_inst : FD1 port map( D => n5014, CP => CLK_I, Q => 
                           n_1323, QN => n4235);
   KEY_EXPAN0_reg_39_6_inst : FD1 port map( D => n5013, CP => CLK_I, Q => 
                           n_1324, QN => n4222);
   KEY_EXPAN0_reg_38_6_inst : FD1 port map( D => n5012, CP => CLK_I, Q => 
                           n_1325, QN => n4221);
   KEY_EXPAN0_reg_37_6_inst : FD1 port map( D => n5011, CP => CLK_I, Q => 
                           n_1326, QN => n4224);
   KEY_EXPAN0_reg_36_6_inst : FD1 port map( D => n5010, CP => CLK_I, Q => 
                           n_1327, QN => n4223);
   KEY_EXPAN0_reg_35_6_inst : FD1 port map( D => n5009, CP => CLK_I, Q => 
                           n_1328, QN => n4226);
   KEY_EXPAN0_reg_34_6_inst : FD1 port map( D => n5008, CP => CLK_I, Q => 
                           n_1329, QN => n4225);
   KEY_EXPAN0_reg_33_6_inst : FD1 port map( D => n5007, CP => CLK_I, Q => 
                           n_1330, QN => n4228);
   KEY_EXPAN0_reg_32_6_inst : FD1 port map( D => n5006, CP => CLK_I, Q => 
                           n_1331, QN => n4227);
   KEY_EXPAN0_reg_31_6_inst : FD1 port map( D => n5005, CP => CLK_I, Q => 
                           n_1332, QN => n4278);
   KEY_EXPAN0_reg_30_6_inst : FD1 port map( D => n5004, CP => CLK_I, Q => 
                           n_1333, QN => n4277);
   KEY_EXPAN0_reg_29_6_inst : FD1 port map( D => n5003, CP => CLK_I, Q => 
                           n_1334, QN => n4280);
   KEY_EXPAN0_reg_28_6_inst : FD1 port map( D => n5002, CP => CLK_I, Q => 
                           n_1335, QN => n4279);
   KEY_EXPAN0_reg_27_6_inst : FD1 port map( D => n5001, CP => CLK_I, Q => 
                           n_1336, QN => n4282);
   KEY_EXPAN0_reg_26_6_inst : FD1 port map( D => n5000, CP => CLK_I, Q => 
                           n_1337, QN => n4281);
   KEY_EXPAN0_reg_25_6_inst : FD1 port map( D => n4999, CP => CLK_I, Q => 
                           n_1338, QN => n4284);
   KEY_EXPAN0_reg_24_6_inst : FD1 port map( D => n4998, CP => CLK_I, Q => 
                           n_1339, QN => n4283);
   KEY_EXPAN0_reg_23_6_inst : FD1 port map( D => n4997, CP => CLK_I, Q => 
                           n_1340, QN => n4270);
   KEY_EXPAN0_reg_22_6_inst : FD1 port map( D => n4996, CP => CLK_I, Q => 
                           n_1341, QN => n4269);
   KEY_EXPAN0_reg_21_6_inst : FD1 port map( D => n4995, CP => CLK_I, Q => 
                           n_1342, QN => n4272);
   KEY_EXPAN0_reg_20_6_inst : FD1 port map( D => n4994, CP => CLK_I, Q => 
                           n_1343, QN => n4271);
   KEY_EXPAN0_reg_19_6_inst : FD1 port map( D => n4993, CP => CLK_I, Q => 
                           n_1344, QN => n4274);
   KEY_EXPAN0_reg_18_6_inst : FD1 port map( D => n4992, CP => CLK_I, Q => 
                           n_1345, QN => n4273);
   KEY_EXPAN0_reg_17_6_inst : FD1 port map( D => n4991, CP => CLK_I, Q => 
                           n_1346, QN => n4276);
   KEY_EXPAN0_reg_16_6_inst : FD1 port map( D => n4990, CP => CLK_I, Q => 
                           n_1347, QN => n4275);
   KEY_EXPAN0_reg_15_6_inst : FD1 port map( D => n4989, CP => CLK_I, Q => 
                           n_1348, QN => n4262);
   KEY_EXPAN0_reg_14_6_inst : FD1 port map( D => n4988, CP => CLK_I, Q => 
                           n_1349, QN => n4261);
   KEY_EXPAN0_reg_13_6_inst : FD1 port map( D => n4987, CP => CLK_I, Q => 
                           n_1350, QN => n4264);
   KEY_EXPAN0_reg_12_6_inst : FD1 port map( D => n4986, CP => CLK_I, Q => 
                           n_1351, QN => n4263);
   KEY_EXPAN0_reg_11_6_inst : FD1 port map( D => n4985, CP => CLK_I, Q => 
                           n_1352, QN => n4266);
   KEY_EXPAN0_reg_10_6_inst : FD1 port map( D => n4984, CP => CLK_I, Q => 
                           n_1353, QN => n4265);
   KEY_EXPAN0_reg_9_6_inst : FD1 port map( D => n4983, CP => CLK_I, Q => n_1354
                           , QN => n4268);
   KEY_EXPAN0_reg_8_6_inst : FD1 port map( D => n4982, CP => CLK_I, Q => n_1355
                           , QN => n4267);
   KEY_EXPAN0_reg_7_6_inst : FD1 port map( D => n4981, CP => CLK_I, Q => n_1356
                           , QN => n4254);
   KEY_EXPAN0_reg_6_6_inst : FD1 port map( D => n4980, CP => CLK_I, Q => n_1357
                           , QN => n4253);
   KEY_EXPAN0_reg_5_6_inst : FD1 port map( D => n4979, CP => CLK_I, Q => n_1358
                           , QN => n4256);
   KEY_EXPAN0_reg_4_6_inst : FD1 port map( D => n4978, CP => CLK_I, Q => n_1359
                           , QN => n4255);
   KEY_EXPAN0_reg_3_6_inst : FD1 port map( D => n4977, CP => CLK_I, Q => n_1360
                           , QN => n4258);
   KEY_EXPAN0_reg_2_6_inst : FD1 port map( D => n4976, CP => CLK_I, Q => n_1361
                           , QN => n4257);
   KEY_EXPAN0_reg_1_6_inst : FD1 port map( D => n4975, CP => CLK_I, Q => n_1362
                           , QN => n4260);
   KEY_EXPAN0_reg_0_6_inst : FD1 port map( D => n4974, CP => CLK_I, Q => n_1363
                           , QN => n4259);
   v_KEY_COL_OUT0_reg_6_inst : FD1 port map( D => n4576, CP => CLK_I, Q => 
                           n4285, QN => n393);
   v_TEMP_VECTOR_reg_30_inst : FD1 port map( D => n6665, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_30_port, QN => n_1364);
   KEY_EXPAN0_reg_63_30_inst : FD1 port map( D => n6573, CP => CLK_I, Q => 
                           n_1365, QN => n4182);
   KEY_EXPAN0_reg_62_30_inst : FD1 port map( D => n6572, CP => CLK_I, Q => 
                           n_1366, QN => n4181);
   KEY_EXPAN0_reg_61_30_inst : FD1 port map( D => n6571, CP => CLK_I, Q => 
                           n_1367, QN => n4184);
   KEY_EXPAN0_reg_60_30_inst : FD1 port map( D => n6570, CP => CLK_I, Q => 
                           n_1368, QN => n4183);
   KEY_EXPAN0_reg_59_30_inst : FD1 port map( D => n6569, CP => CLK_I, Q => 
                           n_1369, QN => n4186);
   KEY_EXPAN0_reg_58_30_inst : FD1 port map( D => n6568, CP => CLK_I, Q => 
                           n_1370, QN => n4185);
   KEY_EXPAN0_reg_57_30_inst : FD1 port map( D => n6567, CP => CLK_I, Q => 
                           n_1371, QN => n4188);
   KEY_EXPAN0_reg_56_30_inst : FD1 port map( D => n6566, CP => CLK_I, Q => 
                           n_1372, QN => n4187);
   KEY_EXPAN0_reg_55_30_inst : FD1 port map( D => n6565, CP => CLK_I, Q => 
                           n_1373, QN => n4174);
   KEY_EXPAN0_reg_54_30_inst : FD1 port map( D => n6564, CP => CLK_I, Q => 
                           n_1374, QN => n4173);
   KEY_EXPAN0_reg_53_30_inst : FD1 port map( D => n6563, CP => CLK_I, Q => 
                           n_1375, QN => n4176);
   KEY_EXPAN0_reg_52_30_inst : FD1 port map( D => n6562, CP => CLK_I, Q => 
                           n_1376, QN => n4175);
   KEY_EXPAN0_reg_51_30_inst : FD1 port map( D => n6561, CP => CLK_I, Q => 
                           n_1377, QN => n4178);
   KEY_EXPAN0_reg_50_30_inst : FD1 port map( D => n6560, CP => CLK_I, Q => 
                           n_1378, QN => n4177);
   KEY_EXPAN0_reg_49_30_inst : FD1 port map( D => n6559, CP => CLK_I, Q => 
                           n_1379, QN => n4180);
   KEY_EXPAN0_reg_48_30_inst : FD1 port map( D => n6558, CP => CLK_I, Q => 
                           n_1380, QN => n4179);
   KEY_EXPAN0_reg_47_30_inst : FD1 port map( D => n6557, CP => CLK_I, Q => 
                           n_1381, QN => n4166);
   KEY_EXPAN0_reg_46_30_inst : FD1 port map( D => n6556, CP => CLK_I, Q => 
                           n_1382, QN => n4165);
   KEY_EXPAN0_reg_45_30_inst : FD1 port map( D => n6555, CP => CLK_I, Q => 
                           n_1383, QN => n4168);
   KEY_EXPAN0_reg_44_30_inst : FD1 port map( D => n6554, CP => CLK_I, Q => 
                           n_1384, QN => n4167);
   KEY_EXPAN0_reg_43_30_inst : FD1 port map( D => n6553, CP => CLK_I, Q => 
                           n_1385, QN => n4170);
   KEY_EXPAN0_reg_42_30_inst : FD1 port map( D => n6552, CP => CLK_I, Q => 
                           n_1386, QN => n4169);
   KEY_EXPAN0_reg_41_30_inst : FD1 port map( D => n6551, CP => CLK_I, Q => 
                           n_1387, QN => n4172);
   KEY_EXPAN0_reg_40_30_inst : FD1 port map( D => n6550, CP => CLK_I, Q => 
                           n_1388, QN => n4171);
   KEY_EXPAN0_reg_39_30_inst : FD1 port map( D => n6549, CP => CLK_I, Q => 
                           n_1389, QN => n4158);
   KEY_EXPAN0_reg_38_30_inst : FD1 port map( D => n6548, CP => CLK_I, Q => 
                           n_1390, QN => n4157);
   KEY_EXPAN0_reg_37_30_inst : FD1 port map( D => n6547, CP => CLK_I, Q => 
                           n_1391, QN => n4160);
   KEY_EXPAN0_reg_36_30_inst : FD1 port map( D => n6546, CP => CLK_I, Q => 
                           n_1392, QN => n4159);
   KEY_EXPAN0_reg_35_30_inst : FD1 port map( D => n6545, CP => CLK_I, Q => 
                           n_1393, QN => n4162);
   KEY_EXPAN0_reg_34_30_inst : FD1 port map( D => n6544, CP => CLK_I, Q => 
                           n_1394, QN => n4161);
   KEY_EXPAN0_reg_33_30_inst : FD1 port map( D => n6543, CP => CLK_I, Q => 
                           n_1395, QN => n4164);
   KEY_EXPAN0_reg_32_30_inst : FD1 port map( D => n6542, CP => CLK_I, Q => 
                           n_1396, QN => n4163);
   KEY_EXPAN0_reg_31_30_inst : FD1 port map( D => n6541, CP => CLK_I, Q => 
                           n_1397, QN => n4214);
   KEY_EXPAN0_reg_30_30_inst : FD1 port map( D => n6540, CP => CLK_I, Q => 
                           n_1398, QN => n4213);
   KEY_EXPAN0_reg_29_30_inst : FD1 port map( D => n6539, CP => CLK_I, Q => 
                           n_1399, QN => n4216);
   KEY_EXPAN0_reg_28_30_inst : FD1 port map( D => n6538, CP => CLK_I, Q => 
                           n_1400, QN => n4215);
   KEY_EXPAN0_reg_27_30_inst : FD1 port map( D => n6537, CP => CLK_I, Q => 
                           n_1401, QN => n4218);
   KEY_EXPAN0_reg_26_30_inst : FD1 port map( D => n6536, CP => CLK_I, Q => 
                           n_1402, QN => n4217);
   KEY_EXPAN0_reg_25_30_inst : FD1 port map( D => n6535, CP => CLK_I, Q => 
                           n_1403, QN => n4220);
   KEY_EXPAN0_reg_24_30_inst : FD1 port map( D => n6534, CP => CLK_I, Q => 
                           n_1404, QN => n4219);
   KEY_EXPAN0_reg_23_30_inst : FD1 port map( D => n6533, CP => CLK_I, Q => 
                           n_1405, QN => n4206);
   KEY_EXPAN0_reg_22_30_inst : FD1 port map( D => n6532, CP => CLK_I, Q => 
                           n_1406, QN => n4205);
   KEY_EXPAN0_reg_21_30_inst : FD1 port map( D => n6531, CP => CLK_I, Q => 
                           n_1407, QN => n4208);
   KEY_EXPAN0_reg_20_30_inst : FD1 port map( D => n6530, CP => CLK_I, Q => 
                           n_1408, QN => n4207);
   KEY_EXPAN0_reg_19_30_inst : FD1 port map( D => n6529, CP => CLK_I, Q => 
                           n_1409, QN => n4210);
   KEY_EXPAN0_reg_18_30_inst : FD1 port map( D => n6528, CP => CLK_I, Q => 
                           n_1410, QN => n4209);
   KEY_EXPAN0_reg_17_30_inst : FD1 port map( D => n6527, CP => CLK_I, Q => 
                           n_1411, QN => n4212);
   KEY_EXPAN0_reg_16_30_inst : FD1 port map( D => n6526, CP => CLK_I, Q => 
                           n_1412, QN => n4211);
   KEY_EXPAN0_reg_15_30_inst : FD1 port map( D => n6525, CP => CLK_I, Q => 
                           n_1413, QN => n4198);
   KEY_EXPAN0_reg_14_30_inst : FD1 port map( D => n6524, CP => CLK_I, Q => 
                           n_1414, QN => n4197);
   KEY_EXPAN0_reg_13_30_inst : FD1 port map( D => n6523, CP => CLK_I, Q => 
                           n_1415, QN => n4200);
   KEY_EXPAN0_reg_12_30_inst : FD1 port map( D => n6522, CP => CLK_I, Q => 
                           n_1416, QN => n4199);
   KEY_EXPAN0_reg_11_30_inst : FD1 port map( D => n6521, CP => CLK_I, Q => 
                           n_1417, QN => n4202);
   KEY_EXPAN0_reg_10_30_inst : FD1 port map( D => n6520, CP => CLK_I, Q => 
                           n_1418, QN => n4201);
   KEY_EXPAN0_reg_9_30_inst : FD1 port map( D => n6519, CP => CLK_I, Q => 
                           n_1419, QN => n4204);
   KEY_EXPAN0_reg_8_30_inst : FD1 port map( D => n6518, CP => CLK_I, Q => 
                           n_1420, QN => n4203);
   KEY_EXPAN0_reg_7_30_inst : FD1 port map( D => n6517, CP => CLK_I, Q => 
                           n_1421, QN => n4190);
   KEY_EXPAN0_reg_6_30_inst : FD1 port map( D => n6516, CP => CLK_I, Q => 
                           n_1422, QN => n4189);
   KEY_EXPAN0_reg_5_30_inst : FD1 port map( D => n6515, CP => CLK_I, Q => 
                           n_1423, QN => n4192);
   KEY_EXPAN0_reg_4_30_inst : FD1 port map( D => n6514, CP => CLK_I, Q => 
                           n_1424, QN => n4191);
   KEY_EXPAN0_reg_3_30_inst : FD1 port map( D => n6513, CP => CLK_I, Q => 
                           n_1425, QN => n4194);
   KEY_EXPAN0_reg_2_30_inst : FD1 port map( D => n6512, CP => CLK_I, Q => 
                           n_1426, QN => n4193);
   KEY_EXPAN0_reg_1_30_inst : FD1 port map( D => n6511, CP => CLK_I, Q => 
                           n_1427, QN => n4196);
   KEY_EXPAN0_reg_0_30_inst : FD1 port map( D => n6510, CP => CLK_I, Q => 
                           n_1428, QN => n4195);
   v_KEY_COL_OUT0_reg_30_inst : FD1 port map( D => n4575, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_30_port, QN => n353);
   v_TEMP_VECTOR_reg_22_inst : FD1 port map( D => n6673, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_22_port, QN => n_1429);
   KEY_EXPAN0_reg_63_22_inst : FD1 port map( D => n6061, CP => CLK_I, Q => 
                           n_1430, QN => n4118);
   KEY_EXPAN0_reg_62_22_inst : FD1 port map( D => n6060, CP => CLK_I, Q => 
                           n_1431, QN => n4117);
   KEY_EXPAN0_reg_61_22_inst : FD1 port map( D => n6059, CP => CLK_I, Q => 
                           n_1432, QN => n4120);
   KEY_EXPAN0_reg_60_22_inst : FD1 port map( D => n6058, CP => CLK_I, Q => 
                           n_1433, QN => n4119);
   KEY_EXPAN0_reg_59_22_inst : FD1 port map( D => n6057, CP => CLK_I, Q => 
                           n_1434, QN => n4122);
   KEY_EXPAN0_reg_58_22_inst : FD1 port map( D => n6056, CP => CLK_I, Q => 
                           n_1435, QN => n4121);
   KEY_EXPAN0_reg_57_22_inst : FD1 port map( D => n6055, CP => CLK_I, Q => 
                           n_1436, QN => n4124);
   KEY_EXPAN0_reg_56_22_inst : FD1 port map( D => n6054, CP => CLK_I, Q => 
                           n_1437, QN => n4123);
   KEY_EXPAN0_reg_55_22_inst : FD1 port map( D => n6053, CP => CLK_I, Q => 
                           n_1438, QN => n4110);
   KEY_EXPAN0_reg_54_22_inst : FD1 port map( D => n6052, CP => CLK_I, Q => 
                           n_1439, QN => n4109);
   KEY_EXPAN0_reg_53_22_inst : FD1 port map( D => n6051, CP => CLK_I, Q => 
                           n_1440, QN => n4112);
   KEY_EXPAN0_reg_52_22_inst : FD1 port map( D => n6050, CP => CLK_I, Q => 
                           n_1441, QN => n4111);
   KEY_EXPAN0_reg_51_22_inst : FD1 port map( D => n6049, CP => CLK_I, Q => 
                           n_1442, QN => n4114);
   KEY_EXPAN0_reg_50_22_inst : FD1 port map( D => n6048, CP => CLK_I, Q => 
                           n_1443, QN => n4113);
   KEY_EXPAN0_reg_49_22_inst : FD1 port map( D => n6047, CP => CLK_I, Q => 
                           n_1444, QN => n4116);
   KEY_EXPAN0_reg_48_22_inst : FD1 port map( D => n6046, CP => CLK_I, Q => 
                           n_1445, QN => n4115);
   KEY_EXPAN0_reg_47_22_inst : FD1 port map( D => n6045, CP => CLK_I, Q => 
                           n_1446, QN => n4102);
   KEY_EXPAN0_reg_46_22_inst : FD1 port map( D => n6044, CP => CLK_I, Q => 
                           n_1447, QN => n4101);
   KEY_EXPAN0_reg_45_22_inst : FD1 port map( D => n6043, CP => CLK_I, Q => 
                           n_1448, QN => n4104);
   KEY_EXPAN0_reg_44_22_inst : FD1 port map( D => n6042, CP => CLK_I, Q => 
                           n_1449, QN => n4103);
   KEY_EXPAN0_reg_43_22_inst : FD1 port map( D => n6041, CP => CLK_I, Q => 
                           n_1450, QN => n4106);
   KEY_EXPAN0_reg_42_22_inst : FD1 port map( D => n6040, CP => CLK_I, Q => 
                           n_1451, QN => n4105);
   KEY_EXPAN0_reg_41_22_inst : FD1 port map( D => n6039, CP => CLK_I, Q => 
                           n_1452, QN => n4108);
   KEY_EXPAN0_reg_40_22_inst : FD1 port map( D => n6038, CP => CLK_I, Q => 
                           n_1453, QN => n4107);
   KEY_EXPAN0_reg_39_22_inst : FD1 port map( D => n6037, CP => CLK_I, Q => 
                           n_1454, QN => n4094);
   KEY_EXPAN0_reg_38_22_inst : FD1 port map( D => n6036, CP => CLK_I, Q => 
                           n_1455, QN => n4093);
   KEY_EXPAN0_reg_37_22_inst : FD1 port map( D => n6035, CP => CLK_I, Q => 
                           n_1456, QN => n4096);
   KEY_EXPAN0_reg_36_22_inst : FD1 port map( D => n6034, CP => CLK_I, Q => 
                           n_1457, QN => n4095);
   KEY_EXPAN0_reg_35_22_inst : FD1 port map( D => n6033, CP => CLK_I, Q => 
                           n_1458, QN => n4098);
   KEY_EXPAN0_reg_34_22_inst : FD1 port map( D => n6032, CP => CLK_I, Q => 
                           n_1459, QN => n4097);
   KEY_EXPAN0_reg_33_22_inst : FD1 port map( D => n6031, CP => CLK_I, Q => 
                           n_1460, QN => n4100);
   KEY_EXPAN0_reg_32_22_inst : FD1 port map( D => n6030, CP => CLK_I, Q => 
                           n_1461, QN => n4099);
   KEY_EXPAN0_reg_31_22_inst : FD1 port map( D => n6029, CP => CLK_I, Q => 
                           n_1462, QN => n4150);
   KEY_EXPAN0_reg_30_22_inst : FD1 port map( D => n6028, CP => CLK_I, Q => 
                           n_1463, QN => n4149);
   KEY_EXPAN0_reg_29_22_inst : FD1 port map( D => n6027, CP => CLK_I, Q => 
                           n_1464, QN => n4152);
   KEY_EXPAN0_reg_28_22_inst : FD1 port map( D => n6026, CP => CLK_I, Q => 
                           n_1465, QN => n4151);
   KEY_EXPAN0_reg_27_22_inst : FD1 port map( D => n6025, CP => CLK_I, Q => 
                           n_1466, QN => n4154);
   KEY_EXPAN0_reg_26_22_inst : FD1 port map( D => n6024, CP => CLK_I, Q => 
                           n_1467, QN => n4153);
   KEY_EXPAN0_reg_25_22_inst : FD1 port map( D => n6023, CP => CLK_I, Q => 
                           n_1468, QN => n4156);
   KEY_EXPAN0_reg_24_22_inst : FD1 port map( D => n6022, CP => CLK_I, Q => 
                           n_1469, QN => n4155);
   KEY_EXPAN0_reg_23_22_inst : FD1 port map( D => n6021, CP => CLK_I, Q => 
                           n_1470, QN => n4142);
   KEY_EXPAN0_reg_22_22_inst : FD1 port map( D => n6020, CP => CLK_I, Q => 
                           n_1471, QN => n4141);
   KEY_EXPAN0_reg_21_22_inst : FD1 port map( D => n6019, CP => CLK_I, Q => 
                           n_1472, QN => n4144);
   KEY_EXPAN0_reg_20_22_inst : FD1 port map( D => n6018, CP => CLK_I, Q => 
                           n_1473, QN => n4143);
   KEY_EXPAN0_reg_19_22_inst : FD1 port map( D => n6017, CP => CLK_I, Q => 
                           n_1474, QN => n4146);
   KEY_EXPAN0_reg_18_22_inst : FD1 port map( D => n6016, CP => CLK_I, Q => 
                           n_1475, QN => n4145);
   KEY_EXPAN0_reg_17_22_inst : FD1 port map( D => n6015, CP => CLK_I, Q => 
                           n_1476, QN => n4148);
   KEY_EXPAN0_reg_16_22_inst : FD1 port map( D => n6014, CP => CLK_I, Q => 
                           n_1477, QN => n4147);
   KEY_EXPAN0_reg_15_22_inst : FD1 port map( D => n6013, CP => CLK_I, Q => 
                           n_1478, QN => n4134);
   KEY_EXPAN0_reg_14_22_inst : FD1 port map( D => n6012, CP => CLK_I, Q => 
                           n_1479, QN => n4133);
   KEY_EXPAN0_reg_13_22_inst : FD1 port map( D => n6011, CP => CLK_I, Q => 
                           n_1480, QN => n4136);
   KEY_EXPAN0_reg_12_22_inst : FD1 port map( D => n6010, CP => CLK_I, Q => 
                           n_1481, QN => n4135);
   KEY_EXPAN0_reg_11_22_inst : FD1 port map( D => n6009, CP => CLK_I, Q => 
                           n_1482, QN => n4138);
   KEY_EXPAN0_reg_10_22_inst : FD1 port map( D => n6008, CP => CLK_I, Q => 
                           n_1483, QN => n4137);
   KEY_EXPAN0_reg_9_22_inst : FD1 port map( D => n6007, CP => CLK_I, Q => 
                           n_1484, QN => n4140);
   KEY_EXPAN0_reg_8_22_inst : FD1 port map( D => n6006, CP => CLK_I, Q => 
                           n_1485, QN => n4139);
   KEY_EXPAN0_reg_7_22_inst : FD1 port map( D => n6005, CP => CLK_I, Q => 
                           n_1486, QN => n4126);
   KEY_EXPAN0_reg_6_22_inst : FD1 port map( D => n6004, CP => CLK_I, Q => 
                           n_1487, QN => n4125);
   KEY_EXPAN0_reg_5_22_inst : FD1 port map( D => n6003, CP => CLK_I, Q => 
                           n_1488, QN => n4128);
   KEY_EXPAN0_reg_4_22_inst : FD1 port map( D => n6002, CP => CLK_I, Q => 
                           n_1489, QN => n4127);
   KEY_EXPAN0_reg_3_22_inst : FD1 port map( D => n6001, CP => CLK_I, Q => 
                           n_1490, QN => n4130);
   KEY_EXPAN0_reg_2_22_inst : FD1 port map( D => n6000, CP => CLK_I, Q => 
                           n_1491, QN => n4129);
   KEY_EXPAN0_reg_1_22_inst : FD1 port map( D => n5999, CP => CLK_I, Q => 
                           n_1492, QN => n4132);
   KEY_EXPAN0_reg_0_22_inst : FD1 port map( D => n5998, CP => CLK_I, Q => 
                           n_1493, QN => n4131);
   v_KEY_COL_OUT0_reg_22_inst : FD1 port map( D => n4574, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_22_port, QN => n352);
   v_TEMP_VECTOR_reg_14_inst : FD1 port map( D => n6681, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_14_port, QN => n_1494);
   KEY_EXPAN0_reg_63_14_inst : FD1 port map( D => n5549, CP => CLK_I, Q => 
                           n_1495, QN => n4054);
   KEY_EXPAN0_reg_62_14_inst : FD1 port map( D => n5548, CP => CLK_I, Q => 
                           n_1496, QN => n4053);
   KEY_EXPAN0_reg_61_14_inst : FD1 port map( D => n5547, CP => CLK_I, Q => 
                           n_1497, QN => n4056);
   KEY_EXPAN0_reg_60_14_inst : FD1 port map( D => n5546, CP => CLK_I, Q => 
                           n_1498, QN => n4055);
   KEY_EXPAN0_reg_59_14_inst : FD1 port map( D => n5545, CP => CLK_I, Q => 
                           n_1499, QN => n4058);
   KEY_EXPAN0_reg_58_14_inst : FD1 port map( D => n5544, CP => CLK_I, Q => 
                           n_1500, QN => n4057);
   KEY_EXPAN0_reg_57_14_inst : FD1 port map( D => n5543, CP => CLK_I, Q => 
                           n_1501, QN => n4060);
   KEY_EXPAN0_reg_56_14_inst : FD1 port map( D => n5542, CP => CLK_I, Q => 
                           n_1502, QN => n4059);
   KEY_EXPAN0_reg_55_14_inst : FD1 port map( D => n5541, CP => CLK_I, Q => 
                           n_1503, QN => n4046);
   KEY_EXPAN0_reg_54_14_inst : FD1 port map( D => n5540, CP => CLK_I, Q => 
                           n_1504, QN => n4045);
   KEY_EXPAN0_reg_53_14_inst : FD1 port map( D => n5539, CP => CLK_I, Q => 
                           n_1505, QN => n4048);
   KEY_EXPAN0_reg_52_14_inst : FD1 port map( D => n5538, CP => CLK_I, Q => 
                           n_1506, QN => n4047);
   KEY_EXPAN0_reg_51_14_inst : FD1 port map( D => n5537, CP => CLK_I, Q => 
                           n_1507, QN => n4050);
   KEY_EXPAN0_reg_50_14_inst : FD1 port map( D => n5536, CP => CLK_I, Q => 
                           n_1508, QN => n4049);
   KEY_EXPAN0_reg_49_14_inst : FD1 port map( D => n5535, CP => CLK_I, Q => 
                           n_1509, QN => n4052);
   KEY_EXPAN0_reg_48_14_inst : FD1 port map( D => n5534, CP => CLK_I, Q => 
                           n_1510, QN => n4051);
   KEY_EXPAN0_reg_47_14_inst : FD1 port map( D => n5533, CP => CLK_I, Q => 
                           n_1511, QN => n4038);
   KEY_EXPAN0_reg_46_14_inst : FD1 port map( D => n5532, CP => CLK_I, Q => 
                           n_1512, QN => n4037);
   KEY_EXPAN0_reg_45_14_inst : FD1 port map( D => n5531, CP => CLK_I, Q => 
                           n_1513, QN => n4040);
   KEY_EXPAN0_reg_44_14_inst : FD1 port map( D => n5530, CP => CLK_I, Q => 
                           n_1514, QN => n4039);
   KEY_EXPAN0_reg_43_14_inst : FD1 port map( D => n5529, CP => CLK_I, Q => 
                           n_1515, QN => n4042);
   KEY_EXPAN0_reg_42_14_inst : FD1 port map( D => n5528, CP => CLK_I, Q => 
                           n_1516, QN => n4041);
   KEY_EXPAN0_reg_41_14_inst : FD1 port map( D => n5527, CP => CLK_I, Q => 
                           n_1517, QN => n4044);
   KEY_EXPAN0_reg_40_14_inst : FD1 port map( D => n5526, CP => CLK_I, Q => 
                           n_1518, QN => n4043);
   KEY_EXPAN0_reg_39_14_inst : FD1 port map( D => n5525, CP => CLK_I, Q => 
                           n_1519, QN => n4030);
   KEY_EXPAN0_reg_38_14_inst : FD1 port map( D => n5524, CP => CLK_I, Q => 
                           n_1520, QN => n4029);
   KEY_EXPAN0_reg_37_14_inst : FD1 port map( D => n5523, CP => CLK_I, Q => 
                           n_1521, QN => n4032);
   KEY_EXPAN0_reg_36_14_inst : FD1 port map( D => n5522, CP => CLK_I, Q => 
                           n_1522, QN => n4031);
   KEY_EXPAN0_reg_35_14_inst : FD1 port map( D => n5521, CP => CLK_I, Q => 
                           n_1523, QN => n4034);
   KEY_EXPAN0_reg_34_14_inst : FD1 port map( D => n5520, CP => CLK_I, Q => 
                           n_1524, QN => n4033);
   KEY_EXPAN0_reg_33_14_inst : FD1 port map( D => n5519, CP => CLK_I, Q => 
                           n_1525, QN => n4036);
   KEY_EXPAN0_reg_32_14_inst : FD1 port map( D => n5518, CP => CLK_I, Q => 
                           n_1526, QN => n4035);
   KEY_EXPAN0_reg_31_14_inst : FD1 port map( D => n5517, CP => CLK_I, Q => 
                           n_1527, QN => n4086);
   KEY_EXPAN0_reg_30_14_inst : FD1 port map( D => n5516, CP => CLK_I, Q => 
                           n_1528, QN => n4085);
   KEY_EXPAN0_reg_29_14_inst : FD1 port map( D => n5515, CP => CLK_I, Q => 
                           n_1529, QN => n4088);
   KEY_EXPAN0_reg_28_14_inst : FD1 port map( D => n5514, CP => CLK_I, Q => 
                           n_1530, QN => n4087);
   KEY_EXPAN0_reg_27_14_inst : FD1 port map( D => n5513, CP => CLK_I, Q => 
                           n_1531, QN => n4090);
   KEY_EXPAN0_reg_26_14_inst : FD1 port map( D => n5512, CP => CLK_I, Q => 
                           n_1532, QN => n4089);
   KEY_EXPAN0_reg_25_14_inst : FD1 port map( D => n5511, CP => CLK_I, Q => 
                           n_1533, QN => n4092);
   KEY_EXPAN0_reg_24_14_inst : FD1 port map( D => n5510, CP => CLK_I, Q => 
                           n_1534, QN => n4091);
   KEY_EXPAN0_reg_23_14_inst : FD1 port map( D => n5509, CP => CLK_I, Q => 
                           n_1535, QN => n4078);
   KEY_EXPAN0_reg_22_14_inst : FD1 port map( D => n5508, CP => CLK_I, Q => 
                           n_1536, QN => n4077);
   KEY_EXPAN0_reg_21_14_inst : FD1 port map( D => n5507, CP => CLK_I, Q => 
                           n_1537, QN => n4080);
   KEY_EXPAN0_reg_20_14_inst : FD1 port map( D => n5506, CP => CLK_I, Q => 
                           n_1538, QN => n4079);
   KEY_EXPAN0_reg_19_14_inst : FD1 port map( D => n5505, CP => CLK_I, Q => 
                           n_1539, QN => n4082);
   KEY_EXPAN0_reg_18_14_inst : FD1 port map( D => n5504, CP => CLK_I, Q => 
                           n_1540, QN => n4081);
   KEY_EXPAN0_reg_17_14_inst : FD1 port map( D => n5503, CP => CLK_I, Q => 
                           n_1541, QN => n4084);
   KEY_EXPAN0_reg_16_14_inst : FD1 port map( D => n5502, CP => CLK_I, Q => 
                           n_1542, QN => n4083);
   KEY_EXPAN0_reg_15_14_inst : FD1 port map( D => n5501, CP => CLK_I, Q => 
                           n_1543, QN => n4070);
   KEY_EXPAN0_reg_14_14_inst : FD1 port map( D => n5500, CP => CLK_I, Q => 
                           n_1544, QN => n4069);
   KEY_EXPAN0_reg_13_14_inst : FD1 port map( D => n5499, CP => CLK_I, Q => 
                           n_1545, QN => n4072);
   KEY_EXPAN0_reg_12_14_inst : FD1 port map( D => n5498, CP => CLK_I, Q => 
                           n_1546, QN => n4071);
   KEY_EXPAN0_reg_11_14_inst : FD1 port map( D => n5497, CP => CLK_I, Q => 
                           n_1547, QN => n4074);
   KEY_EXPAN0_reg_10_14_inst : FD1 port map( D => n5496, CP => CLK_I, Q => 
                           n_1548, QN => n4073);
   KEY_EXPAN0_reg_9_14_inst : FD1 port map( D => n5495, CP => CLK_I, Q => 
                           n_1549, QN => n4076);
   KEY_EXPAN0_reg_8_14_inst : FD1 port map( D => n5494, CP => CLK_I, Q => 
                           n_1550, QN => n4075);
   KEY_EXPAN0_reg_7_14_inst : FD1 port map( D => n5493, CP => CLK_I, Q => 
                           n_1551, QN => n4062);
   KEY_EXPAN0_reg_6_14_inst : FD1 port map( D => n5492, CP => CLK_I, Q => 
                           n_1552, QN => n4061);
   KEY_EXPAN0_reg_5_14_inst : FD1 port map( D => n5491, CP => CLK_I, Q => 
                           n_1553, QN => n4064);
   KEY_EXPAN0_reg_4_14_inst : FD1 port map( D => n5490, CP => CLK_I, Q => 
                           n_1554, QN => n4063);
   KEY_EXPAN0_reg_3_14_inst : FD1 port map( D => n5489, CP => CLK_I, Q => 
                           n_1555, QN => n4066);
   KEY_EXPAN0_reg_2_14_inst : FD1 port map( D => n5488, CP => CLK_I, Q => 
                           n_1556, QN => n4065);
   KEY_EXPAN0_reg_1_14_inst : FD1 port map( D => n5487, CP => CLK_I, Q => 
                           n_1557, QN => n4068);
   KEY_EXPAN0_reg_0_14_inst : FD1 port map( D => n5486, CP => CLK_I, Q => 
                           n_1558, QN => n4067);
   v_KEY_COL_OUT0_reg_14_inst : FD1 port map( D => n4573, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_14_port, QN => n339);
   v_TEMP_VECTOR_reg_5_inst : FD1 port map( D => n6690, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_5_port, QN => n_1559);
   KEY_EXPAN0_reg_63_5_inst : FD1 port map( D => n4973, CP => CLK_I, Q => 
                           n_1560, QN => n3990);
   KEY_EXPAN0_reg_62_5_inst : FD1 port map( D => n4972, CP => CLK_I, Q => 
                           n_1561, QN => n3989);
   KEY_EXPAN0_reg_61_5_inst : FD1 port map( D => n4971, CP => CLK_I, Q => 
                           n_1562, QN => n3992);
   KEY_EXPAN0_reg_60_5_inst : FD1 port map( D => n4970, CP => CLK_I, Q => 
                           n_1563, QN => n3991);
   KEY_EXPAN0_reg_59_5_inst : FD1 port map( D => n4969, CP => CLK_I, Q => 
                           n_1564, QN => n3994);
   KEY_EXPAN0_reg_58_5_inst : FD1 port map( D => n4968, CP => CLK_I, Q => 
                           n_1565, QN => n3993);
   KEY_EXPAN0_reg_57_5_inst : FD1 port map( D => n4967, CP => CLK_I, Q => 
                           n_1566, QN => n3996);
   KEY_EXPAN0_reg_56_5_inst : FD1 port map( D => n4966, CP => CLK_I, Q => 
                           n_1567, QN => n3995);
   KEY_EXPAN0_reg_55_5_inst : FD1 port map( D => n4965, CP => CLK_I, Q => 
                           n_1568, QN => n3982);
   KEY_EXPAN0_reg_54_5_inst : FD1 port map( D => n4964, CP => CLK_I, Q => 
                           n_1569, QN => n3981);
   KEY_EXPAN0_reg_53_5_inst : FD1 port map( D => n4963, CP => CLK_I, Q => 
                           n_1570, QN => n3984);
   KEY_EXPAN0_reg_52_5_inst : FD1 port map( D => n4962, CP => CLK_I, Q => 
                           n_1571, QN => n3983);
   KEY_EXPAN0_reg_51_5_inst : FD1 port map( D => n4961, CP => CLK_I, Q => 
                           n_1572, QN => n3986);
   KEY_EXPAN0_reg_50_5_inst : FD1 port map( D => n4960, CP => CLK_I, Q => 
                           n_1573, QN => n3985);
   KEY_EXPAN0_reg_49_5_inst : FD1 port map( D => n4959, CP => CLK_I, Q => 
                           n_1574, QN => n3988);
   KEY_EXPAN0_reg_48_5_inst : FD1 port map( D => n4958, CP => CLK_I, Q => 
                           n_1575, QN => n3987);
   KEY_EXPAN0_reg_47_5_inst : FD1 port map( D => n4957, CP => CLK_I, Q => 
                           n_1576, QN => n3974);
   KEY_EXPAN0_reg_46_5_inst : FD1 port map( D => n4956, CP => CLK_I, Q => 
                           n_1577, QN => n3973);
   KEY_EXPAN0_reg_45_5_inst : FD1 port map( D => n4955, CP => CLK_I, Q => 
                           n_1578, QN => n3976);
   KEY_EXPAN0_reg_44_5_inst : FD1 port map( D => n4954, CP => CLK_I, Q => 
                           n_1579, QN => n3975);
   KEY_EXPAN0_reg_43_5_inst : FD1 port map( D => n4953, CP => CLK_I, Q => 
                           n_1580, QN => n3978);
   KEY_EXPAN0_reg_42_5_inst : FD1 port map( D => n4952, CP => CLK_I, Q => 
                           n_1581, QN => n3977);
   KEY_EXPAN0_reg_41_5_inst : FD1 port map( D => n4951, CP => CLK_I, Q => 
                           n_1582, QN => n3980);
   KEY_EXPAN0_reg_40_5_inst : FD1 port map( D => n4950, CP => CLK_I, Q => 
                           n_1583, QN => n3979);
   KEY_EXPAN0_reg_39_5_inst : FD1 port map( D => n4949, CP => CLK_I, Q => 
                           n_1584, QN => n3966);
   KEY_EXPAN0_reg_38_5_inst : FD1 port map( D => n4948, CP => CLK_I, Q => 
                           n_1585, QN => n3965);
   KEY_EXPAN0_reg_37_5_inst : FD1 port map( D => n4947, CP => CLK_I, Q => 
                           n_1586, QN => n3968);
   KEY_EXPAN0_reg_36_5_inst : FD1 port map( D => n4946, CP => CLK_I, Q => 
                           n_1587, QN => n3967);
   KEY_EXPAN0_reg_35_5_inst : FD1 port map( D => n4945, CP => CLK_I, Q => 
                           n_1588, QN => n3970);
   KEY_EXPAN0_reg_34_5_inst : FD1 port map( D => n4944, CP => CLK_I, Q => 
                           n_1589, QN => n3969);
   KEY_EXPAN0_reg_33_5_inst : FD1 port map( D => n4943, CP => CLK_I, Q => 
                           n_1590, QN => n3972);
   KEY_EXPAN0_reg_32_5_inst : FD1 port map( D => n4942, CP => CLK_I, Q => 
                           n_1591, QN => n3971);
   KEY_EXPAN0_reg_31_5_inst : FD1 port map( D => n4941, CP => CLK_I, Q => 
                           n_1592, QN => n4022);
   KEY_EXPAN0_reg_30_5_inst : FD1 port map( D => n4940, CP => CLK_I, Q => 
                           n_1593, QN => n4021);
   KEY_EXPAN0_reg_29_5_inst : FD1 port map( D => n4939, CP => CLK_I, Q => 
                           n_1594, QN => n4024);
   KEY_EXPAN0_reg_28_5_inst : FD1 port map( D => n4938, CP => CLK_I, Q => 
                           n_1595, QN => n4023);
   KEY_EXPAN0_reg_27_5_inst : FD1 port map( D => n4937, CP => CLK_I, Q => 
                           n_1596, QN => n4026);
   KEY_EXPAN0_reg_26_5_inst : FD1 port map( D => n4936, CP => CLK_I, Q => 
                           n_1597, QN => n4025);
   KEY_EXPAN0_reg_25_5_inst : FD1 port map( D => n4935, CP => CLK_I, Q => 
                           n_1598, QN => n4028);
   KEY_EXPAN0_reg_24_5_inst : FD1 port map( D => n4934, CP => CLK_I, Q => 
                           n_1599, QN => n4027);
   KEY_EXPAN0_reg_23_5_inst : FD1 port map( D => n4933, CP => CLK_I, Q => 
                           n_1600, QN => n4014);
   KEY_EXPAN0_reg_22_5_inst : FD1 port map( D => n4932, CP => CLK_I, Q => 
                           n_1601, QN => n4013);
   KEY_EXPAN0_reg_21_5_inst : FD1 port map( D => n4931, CP => CLK_I, Q => 
                           n_1602, QN => n4016);
   KEY_EXPAN0_reg_20_5_inst : FD1 port map( D => n4930, CP => CLK_I, Q => 
                           n_1603, QN => n4015);
   KEY_EXPAN0_reg_19_5_inst : FD1 port map( D => n4929, CP => CLK_I, Q => 
                           n_1604, QN => n4018);
   KEY_EXPAN0_reg_18_5_inst : FD1 port map( D => n4928, CP => CLK_I, Q => 
                           n_1605, QN => n4017);
   KEY_EXPAN0_reg_17_5_inst : FD1 port map( D => n4927, CP => CLK_I, Q => 
                           n_1606, QN => n4020);
   KEY_EXPAN0_reg_16_5_inst : FD1 port map( D => n4926, CP => CLK_I, Q => 
                           n_1607, QN => n4019);
   KEY_EXPAN0_reg_15_5_inst : FD1 port map( D => n4925, CP => CLK_I, Q => 
                           n_1608, QN => n4006);
   KEY_EXPAN0_reg_14_5_inst : FD1 port map( D => n4924, CP => CLK_I, Q => 
                           n_1609, QN => n4005);
   KEY_EXPAN0_reg_13_5_inst : FD1 port map( D => n4923, CP => CLK_I, Q => 
                           n_1610, QN => n4008);
   KEY_EXPAN0_reg_12_5_inst : FD1 port map( D => n4922, CP => CLK_I, Q => 
                           n_1611, QN => n4007);
   KEY_EXPAN0_reg_11_5_inst : FD1 port map( D => n4921, CP => CLK_I, Q => 
                           n_1612, QN => n4010);
   KEY_EXPAN0_reg_10_5_inst : FD1 port map( D => n4920, CP => CLK_I, Q => 
                           n_1613, QN => n4009);
   KEY_EXPAN0_reg_9_5_inst : FD1 port map( D => n4919, CP => CLK_I, Q => n_1614
                           , QN => n4012);
   KEY_EXPAN0_reg_8_5_inst : FD1 port map( D => n4918, CP => CLK_I, Q => n_1615
                           , QN => n4011);
   KEY_EXPAN0_reg_7_5_inst : FD1 port map( D => n4917, CP => CLK_I, Q => n_1616
                           , QN => n3998);
   KEY_EXPAN0_reg_6_5_inst : FD1 port map( D => n4916, CP => CLK_I, Q => n_1617
                           , QN => n3997);
   KEY_EXPAN0_reg_5_5_inst : FD1 port map( D => n4915, CP => CLK_I, Q => n_1618
                           , QN => n4000);
   KEY_EXPAN0_reg_4_5_inst : FD1 port map( D => n4914, CP => CLK_I, Q => n_1619
                           , QN => n3999);
   KEY_EXPAN0_reg_3_5_inst : FD1 port map( D => n4913, CP => CLK_I, Q => n_1620
                           , QN => n4002);
   KEY_EXPAN0_reg_2_5_inst : FD1 port map( D => n4912, CP => CLK_I, Q => n_1621
                           , QN => n4001);
   KEY_EXPAN0_reg_1_5_inst : FD1 port map( D => n4911, CP => CLK_I, Q => n_1622
                           , QN => n4004);
   KEY_EXPAN0_reg_0_5_inst : FD1 port map( D => n4910, CP => CLK_I, Q => n_1623
                           , QN => n4003);
   v_KEY_COL_OUT0_reg_5_inst : FD1 port map( D => n4572, CP => CLK_I, Q => 
                           n_1624, QN => n382);
   v_TEMP_VECTOR_reg_29_inst : FD1 port map( D => n6666, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_29_port, QN => n_1625);
   KEY_EXPAN0_reg_63_29_inst : FD1 port map( D => n6509, CP => CLK_I, Q => 
                           n_1626, QN => n3926);
   KEY_EXPAN0_reg_62_29_inst : FD1 port map( D => n6508, CP => CLK_I, Q => 
                           n_1627, QN => n3925);
   KEY_EXPAN0_reg_61_29_inst : FD1 port map( D => n6507, CP => CLK_I, Q => 
                           n_1628, QN => n3928);
   KEY_EXPAN0_reg_60_29_inst : FD1 port map( D => n6506, CP => CLK_I, Q => 
                           n_1629, QN => n3927);
   KEY_EXPAN0_reg_59_29_inst : FD1 port map( D => n6505, CP => CLK_I, Q => 
                           n_1630, QN => n3930);
   KEY_EXPAN0_reg_58_29_inst : FD1 port map( D => n6504, CP => CLK_I, Q => 
                           n_1631, QN => n3929);
   KEY_EXPAN0_reg_57_29_inst : FD1 port map( D => n6503, CP => CLK_I, Q => 
                           n_1632, QN => n3932);
   KEY_EXPAN0_reg_56_29_inst : FD1 port map( D => n6502, CP => CLK_I, Q => 
                           n_1633, QN => n3931);
   KEY_EXPAN0_reg_55_29_inst : FD1 port map( D => n6501, CP => CLK_I, Q => 
                           n_1634, QN => n3918);
   KEY_EXPAN0_reg_54_29_inst : FD1 port map( D => n6500, CP => CLK_I, Q => 
                           n_1635, QN => n3917);
   KEY_EXPAN0_reg_53_29_inst : FD1 port map( D => n6499, CP => CLK_I, Q => 
                           n_1636, QN => n3920);
   KEY_EXPAN0_reg_52_29_inst : FD1 port map( D => n6498, CP => CLK_I, Q => 
                           n_1637, QN => n3919);
   KEY_EXPAN0_reg_51_29_inst : FD1 port map( D => n6497, CP => CLK_I, Q => 
                           n_1638, QN => n3922);
   KEY_EXPAN0_reg_50_29_inst : FD1 port map( D => n6496, CP => CLK_I, Q => 
                           n_1639, QN => n3921);
   KEY_EXPAN0_reg_49_29_inst : FD1 port map( D => n6495, CP => CLK_I, Q => 
                           n_1640, QN => n3924);
   KEY_EXPAN0_reg_48_29_inst : FD1 port map( D => n6494, CP => CLK_I, Q => 
                           n_1641, QN => n3923);
   KEY_EXPAN0_reg_47_29_inst : FD1 port map( D => n6493, CP => CLK_I, Q => 
                           n_1642, QN => n3910);
   KEY_EXPAN0_reg_46_29_inst : FD1 port map( D => n6492, CP => CLK_I, Q => 
                           n_1643, QN => n3909);
   KEY_EXPAN0_reg_45_29_inst : FD1 port map( D => n6491, CP => CLK_I, Q => 
                           n_1644, QN => n3912);
   KEY_EXPAN0_reg_44_29_inst : FD1 port map( D => n6490, CP => CLK_I, Q => 
                           n_1645, QN => n3911);
   KEY_EXPAN0_reg_43_29_inst : FD1 port map( D => n6489, CP => CLK_I, Q => 
                           n_1646, QN => n3914);
   KEY_EXPAN0_reg_42_29_inst : FD1 port map( D => n6488, CP => CLK_I, Q => 
                           n_1647, QN => n3913);
   KEY_EXPAN0_reg_41_29_inst : FD1 port map( D => n6487, CP => CLK_I, Q => 
                           n_1648, QN => n3916);
   KEY_EXPAN0_reg_40_29_inst : FD1 port map( D => n6486, CP => CLK_I, Q => 
                           n_1649, QN => n3915);
   KEY_EXPAN0_reg_39_29_inst : FD1 port map( D => n6485, CP => CLK_I, Q => 
                           n_1650, QN => n3902);
   KEY_EXPAN0_reg_38_29_inst : FD1 port map( D => n6484, CP => CLK_I, Q => 
                           n_1651, QN => n3901);
   KEY_EXPAN0_reg_37_29_inst : FD1 port map( D => n6483, CP => CLK_I, Q => 
                           n_1652, QN => n3904);
   KEY_EXPAN0_reg_36_29_inst : FD1 port map( D => n6482, CP => CLK_I, Q => 
                           n_1653, QN => n3903);
   KEY_EXPAN0_reg_35_29_inst : FD1 port map( D => n6481, CP => CLK_I, Q => 
                           n_1654, QN => n3906);
   KEY_EXPAN0_reg_34_29_inst : FD1 port map( D => n6480, CP => CLK_I, Q => 
                           n_1655, QN => n3905);
   KEY_EXPAN0_reg_33_29_inst : FD1 port map( D => n6479, CP => CLK_I, Q => 
                           n_1656, QN => n3908);
   KEY_EXPAN0_reg_32_29_inst : FD1 port map( D => n6478, CP => CLK_I, Q => 
                           n_1657, QN => n3907);
   KEY_EXPAN0_reg_31_29_inst : FD1 port map( D => n6477, CP => CLK_I, Q => 
                           n_1658, QN => n3958);
   KEY_EXPAN0_reg_30_29_inst : FD1 port map( D => n6476, CP => CLK_I, Q => 
                           n_1659, QN => n3957);
   KEY_EXPAN0_reg_29_29_inst : FD1 port map( D => n6475, CP => CLK_I, Q => 
                           n_1660, QN => n3960);
   KEY_EXPAN0_reg_28_29_inst : FD1 port map( D => n6474, CP => CLK_I, Q => 
                           n_1661, QN => n3959);
   KEY_EXPAN0_reg_27_29_inst : FD1 port map( D => n6473, CP => CLK_I, Q => 
                           n_1662, QN => n3962);
   KEY_EXPAN0_reg_26_29_inst : FD1 port map( D => n6472, CP => CLK_I, Q => 
                           n_1663, QN => n3961);
   KEY_EXPAN0_reg_25_29_inst : FD1 port map( D => n6471, CP => CLK_I, Q => 
                           n_1664, QN => n3964);
   KEY_EXPAN0_reg_24_29_inst : FD1 port map( D => n6470, CP => CLK_I, Q => 
                           n_1665, QN => n3963);
   KEY_EXPAN0_reg_23_29_inst : FD1 port map( D => n6469, CP => CLK_I, Q => 
                           n_1666, QN => n3950);
   KEY_EXPAN0_reg_22_29_inst : FD1 port map( D => n6468, CP => CLK_I, Q => 
                           n_1667, QN => n3949);
   KEY_EXPAN0_reg_21_29_inst : FD1 port map( D => n6467, CP => CLK_I, Q => 
                           n_1668, QN => n3952);
   KEY_EXPAN0_reg_20_29_inst : FD1 port map( D => n6466, CP => CLK_I, Q => 
                           n_1669, QN => n3951);
   KEY_EXPAN0_reg_19_29_inst : FD1 port map( D => n6465, CP => CLK_I, Q => 
                           n_1670, QN => n3954);
   KEY_EXPAN0_reg_18_29_inst : FD1 port map( D => n6464, CP => CLK_I, Q => 
                           n_1671, QN => n3953);
   KEY_EXPAN0_reg_17_29_inst : FD1 port map( D => n6463, CP => CLK_I, Q => 
                           n_1672, QN => n3956);
   KEY_EXPAN0_reg_16_29_inst : FD1 port map( D => n6462, CP => CLK_I, Q => 
                           n_1673, QN => n3955);
   KEY_EXPAN0_reg_15_29_inst : FD1 port map( D => n6461, CP => CLK_I, Q => 
                           n_1674, QN => n3942);
   KEY_EXPAN0_reg_14_29_inst : FD1 port map( D => n6460, CP => CLK_I, Q => 
                           n_1675, QN => n3941);
   KEY_EXPAN0_reg_13_29_inst : FD1 port map( D => n6459, CP => CLK_I, Q => 
                           n_1676, QN => n3944);
   KEY_EXPAN0_reg_12_29_inst : FD1 port map( D => n6458, CP => CLK_I, Q => 
                           n_1677, QN => n3943);
   KEY_EXPAN0_reg_11_29_inst : FD1 port map( D => n6457, CP => CLK_I, Q => 
                           n_1678, QN => n3946);
   KEY_EXPAN0_reg_10_29_inst : FD1 port map( D => n6456, CP => CLK_I, Q => 
                           n_1679, QN => n3945);
   KEY_EXPAN0_reg_9_29_inst : FD1 port map( D => n6455, CP => CLK_I, Q => 
                           n_1680, QN => n3948);
   KEY_EXPAN0_reg_8_29_inst : FD1 port map( D => n6454, CP => CLK_I, Q => 
                           n_1681, QN => n3947);
   KEY_EXPAN0_reg_7_29_inst : FD1 port map( D => n6453, CP => CLK_I, Q => 
                           n_1682, QN => n3934);
   KEY_EXPAN0_reg_6_29_inst : FD1 port map( D => n6452, CP => CLK_I, Q => 
                           n_1683, QN => n3933);
   KEY_EXPAN0_reg_5_29_inst : FD1 port map( D => n6451, CP => CLK_I, Q => 
                           n_1684, QN => n3936);
   KEY_EXPAN0_reg_4_29_inst : FD1 port map( D => n6450, CP => CLK_I, Q => 
                           n_1685, QN => n3935);
   KEY_EXPAN0_reg_3_29_inst : FD1 port map( D => n6449, CP => CLK_I, Q => 
                           n_1686, QN => n3938);
   KEY_EXPAN0_reg_2_29_inst : FD1 port map( D => n6448, CP => CLK_I, Q => 
                           n_1687, QN => n3937);
   KEY_EXPAN0_reg_1_29_inst : FD1 port map( D => n6447, CP => CLK_I, Q => 
                           n_1688, QN => n3940);
   KEY_EXPAN0_reg_0_29_inst : FD1 port map( D => n6446, CP => CLK_I, Q => 
                           n_1689, QN => n3939);
   v_KEY_COL_OUT0_reg_29_inst : FD1 port map( D => n4571, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_29_port, QN => n392);
   v_TEMP_VECTOR_reg_21_inst : FD1 port map( D => n6674, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_21_port, QN => n_1690);
   KEY_EXPAN0_reg_63_21_inst : FD1 port map( D => n5997, CP => CLK_I, Q => 
                           n_1691, QN => n3862);
   KEY_EXPAN0_reg_62_21_inst : FD1 port map( D => n5996, CP => CLK_I, Q => 
                           n_1692, QN => n3861);
   KEY_EXPAN0_reg_61_21_inst : FD1 port map( D => n5995, CP => CLK_I, Q => 
                           n_1693, QN => n3864);
   KEY_EXPAN0_reg_60_21_inst : FD1 port map( D => n5994, CP => CLK_I, Q => 
                           n_1694, QN => n3863);
   KEY_EXPAN0_reg_59_21_inst : FD1 port map( D => n5993, CP => CLK_I, Q => 
                           n_1695, QN => n3866);
   KEY_EXPAN0_reg_58_21_inst : FD1 port map( D => n5992, CP => CLK_I, Q => 
                           n_1696, QN => n3865);
   KEY_EXPAN0_reg_57_21_inst : FD1 port map( D => n5991, CP => CLK_I, Q => 
                           n_1697, QN => n3868);
   KEY_EXPAN0_reg_56_21_inst : FD1 port map( D => n5990, CP => CLK_I, Q => 
                           n_1698, QN => n3867);
   KEY_EXPAN0_reg_55_21_inst : FD1 port map( D => n5989, CP => CLK_I, Q => 
                           n_1699, QN => n3854);
   KEY_EXPAN0_reg_54_21_inst : FD1 port map( D => n5988, CP => CLK_I, Q => 
                           n_1700, QN => n3853);
   KEY_EXPAN0_reg_53_21_inst : FD1 port map( D => n5987, CP => CLK_I, Q => 
                           n_1701, QN => n3856);
   KEY_EXPAN0_reg_52_21_inst : FD1 port map( D => n5986, CP => CLK_I, Q => 
                           n_1702, QN => n3855);
   KEY_EXPAN0_reg_51_21_inst : FD1 port map( D => n5985, CP => CLK_I, Q => 
                           n_1703, QN => n3858);
   KEY_EXPAN0_reg_50_21_inst : FD1 port map( D => n5984, CP => CLK_I, Q => 
                           n_1704, QN => n3857);
   KEY_EXPAN0_reg_49_21_inst : FD1 port map( D => n5983, CP => CLK_I, Q => 
                           n_1705, QN => n3860);
   KEY_EXPAN0_reg_48_21_inst : FD1 port map( D => n5982, CP => CLK_I, Q => 
                           n_1706, QN => n3859);
   KEY_EXPAN0_reg_47_21_inst : FD1 port map( D => n5981, CP => CLK_I, Q => 
                           n_1707, QN => n3846);
   KEY_EXPAN0_reg_46_21_inst : FD1 port map( D => n5980, CP => CLK_I, Q => 
                           n_1708, QN => n3845);
   KEY_EXPAN0_reg_45_21_inst : FD1 port map( D => n5979, CP => CLK_I, Q => 
                           n_1709, QN => n3848);
   KEY_EXPAN0_reg_44_21_inst : FD1 port map( D => n5978, CP => CLK_I, Q => 
                           n_1710, QN => n3847);
   KEY_EXPAN0_reg_43_21_inst : FD1 port map( D => n5977, CP => CLK_I, Q => 
                           n_1711, QN => n3850);
   KEY_EXPAN0_reg_42_21_inst : FD1 port map( D => n5976, CP => CLK_I, Q => 
                           n_1712, QN => n3849);
   KEY_EXPAN0_reg_41_21_inst : FD1 port map( D => n5975, CP => CLK_I, Q => 
                           n_1713, QN => n3852);
   KEY_EXPAN0_reg_40_21_inst : FD1 port map( D => n5974, CP => CLK_I, Q => 
                           n_1714, QN => n3851);
   KEY_EXPAN0_reg_39_21_inst : FD1 port map( D => n5973, CP => CLK_I, Q => 
                           n_1715, QN => n3838);
   KEY_EXPAN0_reg_38_21_inst : FD1 port map( D => n5972, CP => CLK_I, Q => 
                           n_1716, QN => n3837);
   KEY_EXPAN0_reg_37_21_inst : FD1 port map( D => n5971, CP => CLK_I, Q => 
                           n_1717, QN => n3840);
   KEY_EXPAN0_reg_36_21_inst : FD1 port map( D => n5970, CP => CLK_I, Q => 
                           n_1718, QN => n3839);
   KEY_EXPAN0_reg_35_21_inst : FD1 port map( D => n5969, CP => CLK_I, Q => 
                           n_1719, QN => n3842);
   KEY_EXPAN0_reg_34_21_inst : FD1 port map( D => n5968, CP => CLK_I, Q => 
                           n_1720, QN => n3841);
   KEY_EXPAN0_reg_33_21_inst : FD1 port map( D => n5967, CP => CLK_I, Q => 
                           n_1721, QN => n3844);
   KEY_EXPAN0_reg_32_21_inst : FD1 port map( D => n5966, CP => CLK_I, Q => 
                           n_1722, QN => n3843);
   KEY_EXPAN0_reg_31_21_inst : FD1 port map( D => n5965, CP => CLK_I, Q => 
                           n_1723, QN => n3894);
   KEY_EXPAN0_reg_30_21_inst : FD1 port map( D => n5964, CP => CLK_I, Q => 
                           n_1724, QN => n3893);
   KEY_EXPAN0_reg_29_21_inst : FD1 port map( D => n5963, CP => CLK_I, Q => 
                           n_1725, QN => n3896);
   KEY_EXPAN0_reg_28_21_inst : FD1 port map( D => n5962, CP => CLK_I, Q => 
                           n_1726, QN => n3895);
   KEY_EXPAN0_reg_27_21_inst : FD1 port map( D => n5961, CP => CLK_I, Q => 
                           n_1727, QN => n3898);
   KEY_EXPAN0_reg_26_21_inst : FD1 port map( D => n5960, CP => CLK_I, Q => 
                           n_1728, QN => n3897);
   KEY_EXPAN0_reg_25_21_inst : FD1 port map( D => n5959, CP => CLK_I, Q => 
                           n_1729, QN => n3900);
   KEY_EXPAN0_reg_24_21_inst : FD1 port map( D => n5958, CP => CLK_I, Q => 
                           n_1730, QN => n3899);
   KEY_EXPAN0_reg_23_21_inst : FD1 port map( D => n5957, CP => CLK_I, Q => 
                           n_1731, QN => n3886);
   KEY_EXPAN0_reg_22_21_inst : FD1 port map( D => n5956, CP => CLK_I, Q => 
                           n_1732, QN => n3885);
   KEY_EXPAN0_reg_21_21_inst : FD1 port map( D => n5955, CP => CLK_I, Q => 
                           n_1733, QN => n3888);
   KEY_EXPAN0_reg_20_21_inst : FD1 port map( D => n5954, CP => CLK_I, Q => 
                           n_1734, QN => n3887);
   KEY_EXPAN0_reg_19_21_inst : FD1 port map( D => n5953, CP => CLK_I, Q => 
                           n_1735, QN => n3890);
   KEY_EXPAN0_reg_18_21_inst : FD1 port map( D => n5952, CP => CLK_I, Q => 
                           n_1736, QN => n3889);
   KEY_EXPAN0_reg_17_21_inst : FD1 port map( D => n5951, CP => CLK_I, Q => 
                           n_1737, QN => n3892);
   KEY_EXPAN0_reg_16_21_inst : FD1 port map( D => n5950, CP => CLK_I, Q => 
                           n_1738, QN => n3891);
   KEY_EXPAN0_reg_15_21_inst : FD1 port map( D => n5949, CP => CLK_I, Q => 
                           n_1739, QN => n3878);
   KEY_EXPAN0_reg_14_21_inst : FD1 port map( D => n5948, CP => CLK_I, Q => 
                           n_1740, QN => n3877);
   KEY_EXPAN0_reg_13_21_inst : FD1 port map( D => n5947, CP => CLK_I, Q => 
                           n_1741, QN => n3880);
   KEY_EXPAN0_reg_12_21_inst : FD1 port map( D => n5946, CP => CLK_I, Q => 
                           n_1742, QN => n3879);
   KEY_EXPAN0_reg_11_21_inst : FD1 port map( D => n5945, CP => CLK_I, Q => 
                           n_1743, QN => n3882);
   KEY_EXPAN0_reg_10_21_inst : FD1 port map( D => n5944, CP => CLK_I, Q => 
                           n_1744, QN => n3881);
   KEY_EXPAN0_reg_9_21_inst : FD1 port map( D => n5943, CP => CLK_I, Q => 
                           n_1745, QN => n3884);
   KEY_EXPAN0_reg_8_21_inst : FD1 port map( D => n5942, CP => CLK_I, Q => 
                           n_1746, QN => n3883);
   KEY_EXPAN0_reg_7_21_inst : FD1 port map( D => n5941, CP => CLK_I, Q => 
                           n_1747, QN => n3870);
   KEY_EXPAN0_reg_6_21_inst : FD1 port map( D => n5940, CP => CLK_I, Q => 
                           n_1748, QN => n3869);
   KEY_EXPAN0_reg_5_21_inst : FD1 port map( D => n5939, CP => CLK_I, Q => 
                           n_1749, QN => n3872);
   KEY_EXPAN0_reg_4_21_inst : FD1 port map( D => n5938, CP => CLK_I, Q => 
                           n_1750, QN => n3871);
   KEY_EXPAN0_reg_3_21_inst : FD1 port map( D => n5937, CP => CLK_I, Q => 
                           n_1751, QN => n3874);
   KEY_EXPAN0_reg_2_21_inst : FD1 port map( D => n5936, CP => CLK_I, Q => 
                           n_1752, QN => n3873);
   KEY_EXPAN0_reg_1_21_inst : FD1 port map( D => n5935, CP => CLK_I, Q => 
                           n_1753, QN => n3876);
   KEY_EXPAN0_reg_0_21_inst : FD1 port map( D => n5934, CP => CLK_I, Q => 
                           n_1754, QN => n3875);
   v_KEY_COL_OUT0_reg_21_inst : FD1 port map( D => n4570, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_21_port, QN => n351);
   v_TEMP_VECTOR_reg_13_inst : FD1 port map( D => n6682, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_13_port, QN => n_1755);
   KEY_EXPAN0_reg_63_13_inst : FD1 port map( D => n5485, CP => CLK_I, Q => 
                           n_1756, QN => n3798);
   KEY_EXPAN0_reg_62_13_inst : FD1 port map( D => n5484, CP => CLK_I, Q => 
                           n_1757, QN => n3797);
   KEY_EXPAN0_reg_61_13_inst : FD1 port map( D => n5483, CP => CLK_I, Q => 
                           n_1758, QN => n3800);
   KEY_EXPAN0_reg_60_13_inst : FD1 port map( D => n5482, CP => CLK_I, Q => 
                           n_1759, QN => n3799);
   KEY_EXPAN0_reg_59_13_inst : FD1 port map( D => n5481, CP => CLK_I, Q => 
                           n_1760, QN => n3802);
   KEY_EXPAN0_reg_58_13_inst : FD1 port map( D => n5480, CP => CLK_I, Q => 
                           n_1761, QN => n3801);
   KEY_EXPAN0_reg_57_13_inst : FD1 port map( D => n5479, CP => CLK_I, Q => 
                           n_1762, QN => n3804);
   KEY_EXPAN0_reg_56_13_inst : FD1 port map( D => n5478, CP => CLK_I, Q => 
                           n_1763, QN => n3803);
   KEY_EXPAN0_reg_55_13_inst : FD1 port map( D => n5477, CP => CLK_I, Q => 
                           n_1764, QN => n3790);
   KEY_EXPAN0_reg_54_13_inst : FD1 port map( D => n5476, CP => CLK_I, Q => 
                           n_1765, QN => n3789);
   KEY_EXPAN0_reg_53_13_inst : FD1 port map( D => n5475, CP => CLK_I, Q => 
                           n_1766, QN => n3792);
   KEY_EXPAN0_reg_52_13_inst : FD1 port map( D => n5474, CP => CLK_I, Q => 
                           n_1767, QN => n3791);
   KEY_EXPAN0_reg_51_13_inst : FD1 port map( D => n5473, CP => CLK_I, Q => 
                           n_1768, QN => n3794);
   KEY_EXPAN0_reg_50_13_inst : FD1 port map( D => n5472, CP => CLK_I, Q => 
                           n_1769, QN => n3793);
   KEY_EXPAN0_reg_49_13_inst : FD1 port map( D => n5471, CP => CLK_I, Q => 
                           n_1770, QN => n3796);
   KEY_EXPAN0_reg_48_13_inst : FD1 port map( D => n5470, CP => CLK_I, Q => 
                           n_1771, QN => n3795);
   KEY_EXPAN0_reg_47_13_inst : FD1 port map( D => n5469, CP => CLK_I, Q => 
                           n_1772, QN => n3782);
   KEY_EXPAN0_reg_46_13_inst : FD1 port map( D => n5468, CP => CLK_I, Q => 
                           n_1773, QN => n3781);
   KEY_EXPAN0_reg_45_13_inst : FD1 port map( D => n5467, CP => CLK_I, Q => 
                           n_1774, QN => n3784);
   KEY_EXPAN0_reg_44_13_inst : FD1 port map( D => n5466, CP => CLK_I, Q => 
                           n_1775, QN => n3783);
   KEY_EXPAN0_reg_43_13_inst : FD1 port map( D => n5465, CP => CLK_I, Q => 
                           n_1776, QN => n3786);
   KEY_EXPAN0_reg_42_13_inst : FD1 port map( D => n5464, CP => CLK_I, Q => 
                           n_1777, QN => n3785);
   KEY_EXPAN0_reg_41_13_inst : FD1 port map( D => n5463, CP => CLK_I, Q => 
                           n_1778, QN => n3788);
   KEY_EXPAN0_reg_40_13_inst : FD1 port map( D => n5462, CP => CLK_I, Q => 
                           n_1779, QN => n3787);
   KEY_EXPAN0_reg_39_13_inst : FD1 port map( D => n5461, CP => CLK_I, Q => 
                           n_1780, QN => n3774);
   KEY_EXPAN0_reg_38_13_inst : FD1 port map( D => n5460, CP => CLK_I, Q => 
                           n_1781, QN => n3773);
   KEY_EXPAN0_reg_37_13_inst : FD1 port map( D => n5459, CP => CLK_I, Q => 
                           n_1782, QN => n3776);
   KEY_EXPAN0_reg_36_13_inst : FD1 port map( D => n5458, CP => CLK_I, Q => 
                           n_1783, QN => n3775);
   KEY_EXPAN0_reg_35_13_inst : FD1 port map( D => n5457, CP => CLK_I, Q => 
                           n_1784, QN => n3778);
   KEY_EXPAN0_reg_34_13_inst : FD1 port map( D => n5456, CP => CLK_I, Q => 
                           n_1785, QN => n3777);
   KEY_EXPAN0_reg_33_13_inst : FD1 port map( D => n5455, CP => CLK_I, Q => 
                           n_1786, QN => n3780);
   KEY_EXPAN0_reg_32_13_inst : FD1 port map( D => n5454, CP => CLK_I, Q => 
                           n_1787, QN => n3779);
   KEY_EXPAN0_reg_31_13_inst : FD1 port map( D => n5453, CP => CLK_I, Q => 
                           n_1788, QN => n3830);
   KEY_EXPAN0_reg_30_13_inst : FD1 port map( D => n5452, CP => CLK_I, Q => 
                           n_1789, QN => n3829);
   KEY_EXPAN0_reg_29_13_inst : FD1 port map( D => n5451, CP => CLK_I, Q => 
                           n_1790, QN => n3832);
   KEY_EXPAN0_reg_28_13_inst : FD1 port map( D => n5450, CP => CLK_I, Q => 
                           n_1791, QN => n3831);
   KEY_EXPAN0_reg_27_13_inst : FD1 port map( D => n5449, CP => CLK_I, Q => 
                           n_1792, QN => n3834);
   KEY_EXPAN0_reg_26_13_inst : FD1 port map( D => n5448, CP => CLK_I, Q => 
                           n_1793, QN => n3833);
   KEY_EXPAN0_reg_25_13_inst : FD1 port map( D => n5447, CP => CLK_I, Q => 
                           n_1794, QN => n3836);
   KEY_EXPAN0_reg_24_13_inst : FD1 port map( D => n5446, CP => CLK_I, Q => 
                           n_1795, QN => n3835);
   KEY_EXPAN0_reg_23_13_inst : FD1 port map( D => n5445, CP => CLK_I, Q => 
                           n_1796, QN => n3822);
   KEY_EXPAN0_reg_22_13_inst : FD1 port map( D => n5444, CP => CLK_I, Q => 
                           n_1797, QN => n3821);
   KEY_EXPAN0_reg_21_13_inst : FD1 port map( D => n5443, CP => CLK_I, Q => 
                           n_1798, QN => n3824);
   KEY_EXPAN0_reg_20_13_inst : FD1 port map( D => n5442, CP => CLK_I, Q => 
                           n_1799, QN => n3823);
   KEY_EXPAN0_reg_19_13_inst : FD1 port map( D => n5441, CP => CLK_I, Q => 
                           n_1800, QN => n3826);
   KEY_EXPAN0_reg_18_13_inst : FD1 port map( D => n5440, CP => CLK_I, Q => 
                           n_1801, QN => n3825);
   KEY_EXPAN0_reg_17_13_inst : FD1 port map( D => n5439, CP => CLK_I, Q => 
                           n_1802, QN => n3828);
   KEY_EXPAN0_reg_16_13_inst : FD1 port map( D => n5438, CP => CLK_I, Q => 
                           n_1803, QN => n3827);
   KEY_EXPAN0_reg_15_13_inst : FD1 port map( D => n5437, CP => CLK_I, Q => 
                           n_1804, QN => n3814);
   KEY_EXPAN0_reg_14_13_inst : FD1 port map( D => n5436, CP => CLK_I, Q => 
                           n_1805, QN => n3813);
   KEY_EXPAN0_reg_13_13_inst : FD1 port map( D => n5435, CP => CLK_I, Q => 
                           n_1806, QN => n3816);
   KEY_EXPAN0_reg_12_13_inst : FD1 port map( D => n5434, CP => CLK_I, Q => 
                           n_1807, QN => n3815);
   KEY_EXPAN0_reg_11_13_inst : FD1 port map( D => n5433, CP => CLK_I, Q => 
                           n_1808, QN => n3818);
   KEY_EXPAN0_reg_10_13_inst : FD1 port map( D => n5432, CP => CLK_I, Q => 
                           n_1809, QN => n3817);
   KEY_EXPAN0_reg_9_13_inst : FD1 port map( D => n5431, CP => CLK_I, Q => 
                           n_1810, QN => n3820);
   KEY_EXPAN0_reg_8_13_inst : FD1 port map( D => n5430, CP => CLK_I, Q => 
                           n_1811, QN => n3819);
   KEY_EXPAN0_reg_7_13_inst : FD1 port map( D => n5429, CP => CLK_I, Q => 
                           n_1812, QN => n3806);
   KEY_EXPAN0_reg_6_13_inst : FD1 port map( D => n5428, CP => CLK_I, Q => 
                           n_1813, QN => n3805);
   KEY_EXPAN0_reg_5_13_inst : FD1 port map( D => n5427, CP => CLK_I, Q => 
                           n_1814, QN => n3808);
   KEY_EXPAN0_reg_4_13_inst : FD1 port map( D => n5426, CP => CLK_I, Q => 
                           n_1815, QN => n3807);
   KEY_EXPAN0_reg_3_13_inst : FD1 port map( D => n5425, CP => CLK_I, Q => 
                           n_1816, QN => n3810);
   KEY_EXPAN0_reg_2_13_inst : FD1 port map( D => n5424, CP => CLK_I, Q => 
                           n_1817, QN => n3809);
   KEY_EXPAN0_reg_1_13_inst : FD1 port map( D => n5423, CP => CLK_I, Q => 
                           n_1818, QN => n3812);
   KEY_EXPAN0_reg_0_13_inst : FD1 port map( D => n5422, CP => CLK_I, Q => 
                           n_1819, QN => n3811);
   v_KEY_COL_OUT0_reg_13_inst : FD1 port map( D => n4569, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_13_port, QN => n380);
   v_TEMP_VECTOR_reg_4_inst : FD1 port map( D => n6691, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_4_port, QN => n_1820);
   KEY_EXPAN0_reg_63_4_inst : FD1 port map( D => n4909, CP => CLK_I, Q => 
                           n_1821, QN => n3734);
   KEY_EXPAN0_reg_62_4_inst : FD1 port map( D => n4908, CP => CLK_I, Q => 
                           n_1822, QN => n3733);
   KEY_EXPAN0_reg_61_4_inst : FD1 port map( D => n4907, CP => CLK_I, Q => 
                           n_1823, QN => n3736);
   KEY_EXPAN0_reg_60_4_inst : FD1 port map( D => n4906, CP => CLK_I, Q => 
                           n_1824, QN => n3735);
   KEY_EXPAN0_reg_59_4_inst : FD1 port map( D => n4905, CP => CLK_I, Q => 
                           n_1825, QN => n3738);
   KEY_EXPAN0_reg_58_4_inst : FD1 port map( D => n4904, CP => CLK_I, Q => 
                           n_1826, QN => n3737);
   KEY_EXPAN0_reg_57_4_inst : FD1 port map( D => n4903, CP => CLK_I, Q => 
                           n_1827, QN => n3740);
   KEY_EXPAN0_reg_56_4_inst : FD1 port map( D => n4902, CP => CLK_I, Q => 
                           n_1828, QN => n3739);
   KEY_EXPAN0_reg_55_4_inst : FD1 port map( D => n4901, CP => CLK_I, Q => 
                           n_1829, QN => n3726);
   KEY_EXPAN0_reg_54_4_inst : FD1 port map( D => n4900, CP => CLK_I, Q => 
                           n_1830, QN => n3725);
   KEY_EXPAN0_reg_53_4_inst : FD1 port map( D => n4899, CP => CLK_I, Q => 
                           n_1831, QN => n3728);
   KEY_EXPAN0_reg_52_4_inst : FD1 port map( D => n4898, CP => CLK_I, Q => 
                           n_1832, QN => n3727);
   KEY_EXPAN0_reg_51_4_inst : FD1 port map( D => n4897, CP => CLK_I, Q => 
                           n_1833, QN => n3730);
   KEY_EXPAN0_reg_50_4_inst : FD1 port map( D => n4896, CP => CLK_I, Q => 
                           n_1834, QN => n3729);
   KEY_EXPAN0_reg_49_4_inst : FD1 port map( D => n4895, CP => CLK_I, Q => 
                           n_1835, QN => n3732);
   KEY_EXPAN0_reg_48_4_inst : FD1 port map( D => n4894, CP => CLK_I, Q => 
                           n_1836, QN => n3731);
   KEY_EXPAN0_reg_47_4_inst : FD1 port map( D => n4893, CP => CLK_I, Q => 
                           n_1837, QN => n3718);
   KEY_EXPAN0_reg_46_4_inst : FD1 port map( D => n4892, CP => CLK_I, Q => 
                           n_1838, QN => n3717);
   KEY_EXPAN0_reg_45_4_inst : FD1 port map( D => n4891, CP => CLK_I, Q => 
                           n_1839, QN => n3720);
   KEY_EXPAN0_reg_44_4_inst : FD1 port map( D => n4890, CP => CLK_I, Q => 
                           n_1840, QN => n3719);
   KEY_EXPAN0_reg_43_4_inst : FD1 port map( D => n4889, CP => CLK_I, Q => 
                           n_1841, QN => n3722);
   KEY_EXPAN0_reg_42_4_inst : FD1 port map( D => n4888, CP => CLK_I, Q => 
                           n_1842, QN => n3721);
   KEY_EXPAN0_reg_41_4_inst : FD1 port map( D => n4887, CP => CLK_I, Q => 
                           n_1843, QN => n3724);
   KEY_EXPAN0_reg_40_4_inst : FD1 port map( D => n4886, CP => CLK_I, Q => 
                           n_1844, QN => n3723);
   KEY_EXPAN0_reg_39_4_inst : FD1 port map( D => n4885, CP => CLK_I, Q => 
                           n_1845, QN => n3710);
   KEY_EXPAN0_reg_38_4_inst : FD1 port map( D => n4884, CP => CLK_I, Q => 
                           n_1846, QN => n3709);
   KEY_EXPAN0_reg_37_4_inst : FD1 port map( D => n4883, CP => CLK_I, Q => 
                           n_1847, QN => n3712);
   KEY_EXPAN0_reg_36_4_inst : FD1 port map( D => n4882, CP => CLK_I, Q => 
                           n_1848, QN => n3711);
   KEY_EXPAN0_reg_35_4_inst : FD1 port map( D => n4881, CP => CLK_I, Q => 
                           n_1849, QN => n3714);
   KEY_EXPAN0_reg_34_4_inst : FD1 port map( D => n4880, CP => CLK_I, Q => 
                           n_1850, QN => n3713);
   KEY_EXPAN0_reg_33_4_inst : FD1 port map( D => n4879, CP => CLK_I, Q => 
                           n_1851, QN => n3716);
   KEY_EXPAN0_reg_32_4_inst : FD1 port map( D => n4878, CP => CLK_I, Q => 
                           n_1852, QN => n3715);
   KEY_EXPAN0_reg_31_4_inst : FD1 port map( D => n4877, CP => CLK_I, Q => 
                           n_1853, QN => n3766);
   KEY_EXPAN0_reg_30_4_inst : FD1 port map( D => n4876, CP => CLK_I, Q => 
                           n_1854, QN => n3765);
   KEY_EXPAN0_reg_29_4_inst : FD1 port map( D => n4875, CP => CLK_I, Q => 
                           n_1855, QN => n3768);
   KEY_EXPAN0_reg_28_4_inst : FD1 port map( D => n4874, CP => CLK_I, Q => 
                           n_1856, QN => n3767);
   KEY_EXPAN0_reg_27_4_inst : FD1 port map( D => n4873, CP => CLK_I, Q => 
                           n_1857, QN => n3770);
   KEY_EXPAN0_reg_26_4_inst : FD1 port map( D => n4872, CP => CLK_I, Q => 
                           n_1858, QN => n3769);
   KEY_EXPAN0_reg_25_4_inst : FD1 port map( D => n4871, CP => CLK_I, Q => 
                           n_1859, QN => n3772);
   KEY_EXPAN0_reg_24_4_inst : FD1 port map( D => n4870, CP => CLK_I, Q => 
                           n_1860, QN => n3771);
   KEY_EXPAN0_reg_23_4_inst : FD1 port map( D => n4869, CP => CLK_I, Q => 
                           n_1861, QN => n3758);
   KEY_EXPAN0_reg_22_4_inst : FD1 port map( D => n4868, CP => CLK_I, Q => 
                           n_1862, QN => n3757);
   KEY_EXPAN0_reg_21_4_inst : FD1 port map( D => n4867, CP => CLK_I, Q => 
                           n_1863, QN => n3760);
   KEY_EXPAN0_reg_20_4_inst : FD1 port map( D => n4866, CP => CLK_I, Q => 
                           n_1864, QN => n3759);
   KEY_EXPAN0_reg_19_4_inst : FD1 port map( D => n4865, CP => CLK_I, Q => 
                           n_1865, QN => n3762);
   KEY_EXPAN0_reg_18_4_inst : FD1 port map( D => n4864, CP => CLK_I, Q => 
                           n_1866, QN => n3761);
   KEY_EXPAN0_reg_17_4_inst : FD1 port map( D => n4863, CP => CLK_I, Q => 
                           n_1867, QN => n3764);
   KEY_EXPAN0_reg_16_4_inst : FD1 port map( D => n4862, CP => CLK_I, Q => 
                           n_1868, QN => n3763);
   KEY_EXPAN0_reg_15_4_inst : FD1 port map( D => n4861, CP => CLK_I, Q => 
                           n_1869, QN => n3750);
   KEY_EXPAN0_reg_14_4_inst : FD1 port map( D => n4860, CP => CLK_I, Q => 
                           n_1870, QN => n3749);
   KEY_EXPAN0_reg_13_4_inst : FD1 port map( D => n4859, CP => CLK_I, Q => 
                           n_1871, QN => n3752);
   KEY_EXPAN0_reg_12_4_inst : FD1 port map( D => n4858, CP => CLK_I, Q => 
                           n_1872, QN => n3751);
   KEY_EXPAN0_reg_11_4_inst : FD1 port map( D => n4857, CP => CLK_I, Q => 
                           n_1873, QN => n3754);
   KEY_EXPAN0_reg_10_4_inst : FD1 port map( D => n4856, CP => CLK_I, Q => 
                           n_1874, QN => n3753);
   KEY_EXPAN0_reg_9_4_inst : FD1 port map( D => n4855, CP => CLK_I, Q => n_1875
                           , QN => n3756);
   KEY_EXPAN0_reg_8_4_inst : FD1 port map( D => n4854, CP => CLK_I, Q => n_1876
                           , QN => n3755);
   KEY_EXPAN0_reg_7_4_inst : FD1 port map( D => n4853, CP => CLK_I, Q => n_1877
                           , QN => n3742);
   KEY_EXPAN0_reg_6_4_inst : FD1 port map( D => n4852, CP => CLK_I, Q => n_1878
                           , QN => n3741);
   KEY_EXPAN0_reg_5_4_inst : FD1 port map( D => n4851, CP => CLK_I, Q => n_1879
                           , QN => n3744);
   KEY_EXPAN0_reg_4_4_inst : FD1 port map( D => n4850, CP => CLK_I, Q => n_1880
                           , QN => n3743);
   KEY_EXPAN0_reg_3_4_inst : FD1 port map( D => n4849, CP => CLK_I, Q => n_1881
                           , QN => n3746);
   KEY_EXPAN0_reg_2_4_inst : FD1 port map( D => n4848, CP => CLK_I, Q => n_1882
                           , QN => n3745);
   KEY_EXPAN0_reg_1_4_inst : FD1 port map( D => n4847, CP => CLK_I, Q => n_1883
                           , QN => n3748);
   KEY_EXPAN0_reg_0_4_inst : FD1 port map( D => n4846, CP => CLK_I, Q => n_1884
                           , QN => n3747);
   v_KEY_COL_OUT0_reg_4_inst : FD1 port map( D => n4568, CP => CLK_I, Q => 
                           n_1885, QN => n1630);
   v_TEMP_VECTOR_reg_28_inst : FD1 port map( D => n6667, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_28_port, QN => n_1886);
   KEY_EXPAN0_reg_63_28_inst : FD1 port map( D => n6445, CP => CLK_I, Q => 
                           n_1887, QN => n3670);
   KEY_EXPAN0_reg_62_28_inst : FD1 port map( D => n6444, CP => CLK_I, Q => 
                           n_1888, QN => n3669);
   KEY_EXPAN0_reg_61_28_inst : FD1 port map( D => n6443, CP => CLK_I, Q => 
                           n_1889, QN => n3672);
   KEY_EXPAN0_reg_60_28_inst : FD1 port map( D => n6442, CP => CLK_I, Q => 
                           n_1890, QN => n3671);
   KEY_EXPAN0_reg_59_28_inst : FD1 port map( D => n6441, CP => CLK_I, Q => 
                           n_1891, QN => n3674);
   KEY_EXPAN0_reg_58_28_inst : FD1 port map( D => n6440, CP => CLK_I, Q => 
                           n_1892, QN => n3673);
   KEY_EXPAN0_reg_57_28_inst : FD1 port map( D => n6439, CP => CLK_I, Q => 
                           n_1893, QN => n3676);
   KEY_EXPAN0_reg_56_28_inst : FD1 port map( D => n6438, CP => CLK_I, Q => 
                           n_1894, QN => n3675);
   KEY_EXPAN0_reg_55_28_inst : FD1 port map( D => n6437, CP => CLK_I, Q => 
                           n_1895, QN => n3662);
   KEY_EXPAN0_reg_54_28_inst : FD1 port map( D => n6436, CP => CLK_I, Q => 
                           n_1896, QN => n3661);
   KEY_EXPAN0_reg_53_28_inst : FD1 port map( D => n6435, CP => CLK_I, Q => 
                           n_1897, QN => n3664);
   KEY_EXPAN0_reg_52_28_inst : FD1 port map( D => n6434, CP => CLK_I, Q => 
                           n_1898, QN => n3663);
   KEY_EXPAN0_reg_51_28_inst : FD1 port map( D => n6433, CP => CLK_I, Q => 
                           n_1899, QN => n3666);
   KEY_EXPAN0_reg_50_28_inst : FD1 port map( D => n6432, CP => CLK_I, Q => 
                           n_1900, QN => n3665);
   KEY_EXPAN0_reg_49_28_inst : FD1 port map( D => n6431, CP => CLK_I, Q => 
                           n_1901, QN => n3668);
   KEY_EXPAN0_reg_48_28_inst : FD1 port map( D => n6430, CP => CLK_I, Q => 
                           n_1902, QN => n3667);
   KEY_EXPAN0_reg_47_28_inst : FD1 port map( D => n6429, CP => CLK_I, Q => 
                           n_1903, QN => n3654);
   KEY_EXPAN0_reg_46_28_inst : FD1 port map( D => n6428, CP => CLK_I, Q => 
                           n_1904, QN => n3653);
   KEY_EXPAN0_reg_45_28_inst : FD1 port map( D => n6427, CP => CLK_I, Q => 
                           n_1905, QN => n3656);
   KEY_EXPAN0_reg_44_28_inst : FD1 port map( D => n6426, CP => CLK_I, Q => 
                           n_1906, QN => n3655);
   KEY_EXPAN0_reg_43_28_inst : FD1 port map( D => n6425, CP => CLK_I, Q => 
                           n_1907, QN => n3658);
   KEY_EXPAN0_reg_42_28_inst : FD1 port map( D => n6424, CP => CLK_I, Q => 
                           n_1908, QN => n3657);
   KEY_EXPAN0_reg_41_28_inst : FD1 port map( D => n6423, CP => CLK_I, Q => 
                           n_1909, QN => n3660);
   KEY_EXPAN0_reg_40_28_inst : FD1 port map( D => n6422, CP => CLK_I, Q => 
                           n_1910, QN => n3659);
   KEY_EXPAN0_reg_39_28_inst : FD1 port map( D => n6421, CP => CLK_I, Q => 
                           n_1911, QN => n3646);
   KEY_EXPAN0_reg_38_28_inst : FD1 port map( D => n6420, CP => CLK_I, Q => 
                           n_1912, QN => n3645);
   KEY_EXPAN0_reg_37_28_inst : FD1 port map( D => n6419, CP => CLK_I, Q => 
                           n_1913, QN => n3648);
   KEY_EXPAN0_reg_36_28_inst : FD1 port map( D => n6418, CP => CLK_I, Q => 
                           n_1914, QN => n3647);
   KEY_EXPAN0_reg_35_28_inst : FD1 port map( D => n6417, CP => CLK_I, Q => 
                           n_1915, QN => n3650);
   KEY_EXPAN0_reg_34_28_inst : FD1 port map( D => n6416, CP => CLK_I, Q => 
                           n_1916, QN => n3649);
   KEY_EXPAN0_reg_33_28_inst : FD1 port map( D => n6415, CP => CLK_I, Q => 
                           n_1917, QN => n3652);
   KEY_EXPAN0_reg_32_28_inst : FD1 port map( D => n6414, CP => CLK_I, Q => 
                           n_1918, QN => n3651);
   KEY_EXPAN0_reg_31_28_inst : FD1 port map( D => n6413, CP => CLK_I, Q => 
                           n_1919, QN => n3702);
   KEY_EXPAN0_reg_30_28_inst : FD1 port map( D => n6412, CP => CLK_I, Q => 
                           n_1920, QN => n3701);
   KEY_EXPAN0_reg_29_28_inst : FD1 port map( D => n6411, CP => CLK_I, Q => 
                           n_1921, QN => n3704);
   KEY_EXPAN0_reg_28_28_inst : FD1 port map( D => n6410, CP => CLK_I, Q => 
                           n_1922, QN => n3703);
   KEY_EXPAN0_reg_27_28_inst : FD1 port map( D => n6409, CP => CLK_I, Q => 
                           n_1923, QN => n3706);
   KEY_EXPAN0_reg_26_28_inst : FD1 port map( D => n6408, CP => CLK_I, Q => 
                           n_1924, QN => n3705);
   KEY_EXPAN0_reg_25_28_inst : FD1 port map( D => n6407, CP => CLK_I, Q => 
                           n_1925, QN => n3708);
   KEY_EXPAN0_reg_24_28_inst : FD1 port map( D => n6406, CP => CLK_I, Q => 
                           n_1926, QN => n3707);
   KEY_EXPAN0_reg_23_28_inst : FD1 port map( D => n6405, CP => CLK_I, Q => 
                           n_1927, QN => n3694);
   KEY_EXPAN0_reg_22_28_inst : FD1 port map( D => n6404, CP => CLK_I, Q => 
                           n_1928, QN => n3693);
   KEY_EXPAN0_reg_21_28_inst : FD1 port map( D => n6403, CP => CLK_I, Q => 
                           n_1929, QN => n3696);
   KEY_EXPAN0_reg_20_28_inst : FD1 port map( D => n6402, CP => CLK_I, Q => 
                           n_1930, QN => n3695);
   KEY_EXPAN0_reg_19_28_inst : FD1 port map( D => n6401, CP => CLK_I, Q => 
                           n_1931, QN => n3698);
   KEY_EXPAN0_reg_18_28_inst : FD1 port map( D => n6400, CP => CLK_I, Q => 
                           n_1932, QN => n3697);
   KEY_EXPAN0_reg_17_28_inst : FD1 port map( D => n6399, CP => CLK_I, Q => 
                           n_1933, QN => n3700);
   KEY_EXPAN0_reg_16_28_inst : FD1 port map( D => n6398, CP => CLK_I, Q => 
                           n_1934, QN => n3699);
   KEY_EXPAN0_reg_15_28_inst : FD1 port map( D => n6397, CP => CLK_I, Q => 
                           n_1935, QN => n3686);
   KEY_EXPAN0_reg_14_28_inst : FD1 port map( D => n6396, CP => CLK_I, Q => 
                           n_1936, QN => n3685);
   KEY_EXPAN0_reg_13_28_inst : FD1 port map( D => n6395, CP => CLK_I, Q => 
                           n_1937, QN => n3688);
   KEY_EXPAN0_reg_12_28_inst : FD1 port map( D => n6394, CP => CLK_I, Q => 
                           n_1938, QN => n3687);
   KEY_EXPAN0_reg_11_28_inst : FD1 port map( D => n6393, CP => CLK_I, Q => 
                           n_1939, QN => n3690);
   KEY_EXPAN0_reg_10_28_inst : FD1 port map( D => n6392, CP => CLK_I, Q => 
                           n_1940, QN => n3689);
   KEY_EXPAN0_reg_9_28_inst : FD1 port map( D => n6391, CP => CLK_I, Q => 
                           n_1941, QN => n3692);
   KEY_EXPAN0_reg_8_28_inst : FD1 port map( D => n6390, CP => CLK_I, Q => 
                           n_1942, QN => n3691);
   KEY_EXPAN0_reg_7_28_inst : FD1 port map( D => n6389, CP => CLK_I, Q => 
                           n_1943, QN => n3678);
   KEY_EXPAN0_reg_6_28_inst : FD1 port map( D => n6388, CP => CLK_I, Q => 
                           n_1944, QN => n3677);
   KEY_EXPAN0_reg_5_28_inst : FD1 port map( D => n6387, CP => CLK_I, Q => 
                           n_1945, QN => n3680);
   KEY_EXPAN0_reg_4_28_inst : FD1 port map( D => n6386, CP => CLK_I, Q => 
                           n_1946, QN => n3679);
   KEY_EXPAN0_reg_3_28_inst : FD1 port map( D => n6385, CP => CLK_I, Q => 
                           n_1947, QN => n3682);
   KEY_EXPAN0_reg_2_28_inst : FD1 port map( D => n6384, CP => CLK_I, Q => 
                           n_1948, QN => n3681);
   KEY_EXPAN0_reg_1_28_inst : FD1 port map( D => n6383, CP => CLK_I, Q => 
                           n_1949, QN => n3684);
   KEY_EXPAN0_reg_0_28_inst : FD1 port map( D => n6382, CP => CLK_I, Q => 
                           n_1950, QN => n3683);
   v_KEY_COL_OUT0_reg_28_inst : FD1 port map( D => n4567, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_28_port, QN => n1897);
   v_TEMP_VECTOR_reg_20_inst : FD1 port map( D => n6675, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_20_port, QN => n_1951);
   KEY_EXPAN0_reg_63_20_inst : FD1 port map( D => n5933, CP => CLK_I, Q => 
                           n_1952, QN => n3606);
   KEY_EXPAN0_reg_62_20_inst : FD1 port map( D => n5932, CP => CLK_I, Q => 
                           n_1953, QN => n3605);
   KEY_EXPAN0_reg_61_20_inst : FD1 port map( D => n5931, CP => CLK_I, Q => 
                           n_1954, QN => n3608);
   KEY_EXPAN0_reg_60_20_inst : FD1 port map( D => n5930, CP => CLK_I, Q => 
                           n_1955, QN => n3607);
   KEY_EXPAN0_reg_59_20_inst : FD1 port map( D => n5929, CP => CLK_I, Q => 
                           n_1956, QN => n3610);
   KEY_EXPAN0_reg_58_20_inst : FD1 port map( D => n5928, CP => CLK_I, Q => 
                           n_1957, QN => n3609);
   KEY_EXPAN0_reg_57_20_inst : FD1 port map( D => n5927, CP => CLK_I, Q => 
                           n_1958, QN => n3612);
   KEY_EXPAN0_reg_56_20_inst : FD1 port map( D => n5926, CP => CLK_I, Q => 
                           n_1959, QN => n3611);
   KEY_EXPAN0_reg_55_20_inst : FD1 port map( D => n5925, CP => CLK_I, Q => 
                           n_1960, QN => n3598);
   KEY_EXPAN0_reg_54_20_inst : FD1 port map( D => n5924, CP => CLK_I, Q => 
                           n_1961, QN => n3597);
   KEY_EXPAN0_reg_53_20_inst : FD1 port map( D => n5923, CP => CLK_I, Q => 
                           n_1962, QN => n3600);
   KEY_EXPAN0_reg_52_20_inst : FD1 port map( D => n5922, CP => CLK_I, Q => 
                           n_1963, QN => n3599);
   KEY_EXPAN0_reg_51_20_inst : FD1 port map( D => n5921, CP => CLK_I, Q => 
                           n_1964, QN => n3602);
   KEY_EXPAN0_reg_50_20_inst : FD1 port map( D => n5920, CP => CLK_I, Q => 
                           n_1965, QN => n3601);
   KEY_EXPAN0_reg_49_20_inst : FD1 port map( D => n5919, CP => CLK_I, Q => 
                           n_1966, QN => n3604);
   KEY_EXPAN0_reg_48_20_inst : FD1 port map( D => n5918, CP => CLK_I, Q => 
                           n_1967, QN => n3603);
   KEY_EXPAN0_reg_47_20_inst : FD1 port map( D => n5917, CP => CLK_I, Q => 
                           n_1968, QN => n3590);
   KEY_EXPAN0_reg_46_20_inst : FD1 port map( D => n5916, CP => CLK_I, Q => 
                           n_1969, QN => n3589);
   KEY_EXPAN0_reg_45_20_inst : FD1 port map( D => n5915, CP => CLK_I, Q => 
                           n_1970, QN => n3592);
   KEY_EXPAN0_reg_44_20_inst : FD1 port map( D => n5914, CP => CLK_I, Q => 
                           n_1971, QN => n3591);
   KEY_EXPAN0_reg_43_20_inst : FD1 port map( D => n5913, CP => CLK_I, Q => 
                           n_1972, QN => n3594);
   KEY_EXPAN0_reg_42_20_inst : FD1 port map( D => n5912, CP => CLK_I, Q => 
                           n_1973, QN => n3593);
   KEY_EXPAN0_reg_41_20_inst : FD1 port map( D => n5911, CP => CLK_I, Q => 
                           n_1974, QN => n3596);
   KEY_EXPAN0_reg_40_20_inst : FD1 port map( D => n5910, CP => CLK_I, Q => 
                           n_1975, QN => n3595);
   KEY_EXPAN0_reg_39_20_inst : FD1 port map( D => n5909, CP => CLK_I, Q => 
                           n_1976, QN => n3582);
   KEY_EXPAN0_reg_38_20_inst : FD1 port map( D => n5908, CP => CLK_I, Q => 
                           n_1977, QN => n3581);
   KEY_EXPAN0_reg_37_20_inst : FD1 port map( D => n5907, CP => CLK_I, Q => 
                           n_1978, QN => n3584);
   KEY_EXPAN0_reg_36_20_inst : FD1 port map( D => n5906, CP => CLK_I, Q => 
                           n_1979, QN => n3583);
   KEY_EXPAN0_reg_35_20_inst : FD1 port map( D => n5905, CP => CLK_I, Q => 
                           n_1980, QN => n3586);
   KEY_EXPAN0_reg_34_20_inst : FD1 port map( D => n5904, CP => CLK_I, Q => 
                           n_1981, QN => n3585);
   KEY_EXPAN0_reg_33_20_inst : FD1 port map( D => n5903, CP => CLK_I, Q => 
                           n_1982, QN => n3588);
   KEY_EXPAN0_reg_32_20_inst : FD1 port map( D => n5902, CP => CLK_I, Q => 
                           n_1983, QN => n3587);
   KEY_EXPAN0_reg_31_20_inst : FD1 port map( D => n5901, CP => CLK_I, Q => 
                           n_1984, QN => n3638);
   KEY_EXPAN0_reg_30_20_inst : FD1 port map( D => n5900, CP => CLK_I, Q => 
                           n_1985, QN => n3637);
   KEY_EXPAN0_reg_29_20_inst : FD1 port map( D => n5899, CP => CLK_I, Q => 
                           n_1986, QN => n3640);
   KEY_EXPAN0_reg_28_20_inst : FD1 port map( D => n5898, CP => CLK_I, Q => 
                           n_1987, QN => n3639);
   KEY_EXPAN0_reg_27_20_inst : FD1 port map( D => n5897, CP => CLK_I, Q => 
                           n_1988, QN => n3642);
   KEY_EXPAN0_reg_26_20_inst : FD1 port map( D => n5896, CP => CLK_I, Q => 
                           n_1989, QN => n3641);
   KEY_EXPAN0_reg_25_20_inst : FD1 port map( D => n5895, CP => CLK_I, Q => 
                           n_1990, QN => n3644);
   KEY_EXPAN0_reg_24_20_inst : FD1 port map( D => n5894, CP => CLK_I, Q => 
                           n_1991, QN => n3643);
   KEY_EXPAN0_reg_23_20_inst : FD1 port map( D => n5893, CP => CLK_I, Q => 
                           n_1992, QN => n3630);
   KEY_EXPAN0_reg_22_20_inst : FD1 port map( D => n5892, CP => CLK_I, Q => 
                           n_1993, QN => n3629);
   KEY_EXPAN0_reg_21_20_inst : FD1 port map( D => n5891, CP => CLK_I, Q => 
                           n_1994, QN => n3632);
   KEY_EXPAN0_reg_20_20_inst : FD1 port map( D => n5890, CP => CLK_I, Q => 
                           n_1995, QN => n3631);
   KEY_EXPAN0_reg_19_20_inst : FD1 port map( D => n5889, CP => CLK_I, Q => 
                           n_1996, QN => n3634);
   KEY_EXPAN0_reg_18_20_inst : FD1 port map( D => n5888, CP => CLK_I, Q => 
                           n_1997, QN => n3633);
   KEY_EXPAN0_reg_17_20_inst : FD1 port map( D => n5887, CP => CLK_I, Q => 
                           n_1998, QN => n3636);
   KEY_EXPAN0_reg_16_20_inst : FD1 port map( D => n5886, CP => CLK_I, Q => 
                           n_1999, QN => n3635);
   KEY_EXPAN0_reg_15_20_inst : FD1 port map( D => n5885, CP => CLK_I, Q => 
                           n_2000, QN => n3622);
   KEY_EXPAN0_reg_14_20_inst : FD1 port map( D => n5884, CP => CLK_I, Q => 
                           n_2001, QN => n3621);
   KEY_EXPAN0_reg_13_20_inst : FD1 port map( D => n5883, CP => CLK_I, Q => 
                           n_2002, QN => n3624);
   KEY_EXPAN0_reg_12_20_inst : FD1 port map( D => n5882, CP => CLK_I, Q => 
                           n_2003, QN => n3623);
   KEY_EXPAN0_reg_11_20_inst : FD1 port map( D => n5881, CP => CLK_I, Q => 
                           n_2004, QN => n3626);
   KEY_EXPAN0_reg_10_20_inst : FD1 port map( D => n5880, CP => CLK_I, Q => 
                           n_2005, QN => n3625);
   KEY_EXPAN0_reg_9_20_inst : FD1 port map( D => n5879, CP => CLK_I, Q => 
                           n_2006, QN => n3628);
   KEY_EXPAN0_reg_8_20_inst : FD1 port map( D => n5878, CP => CLK_I, Q => 
                           n_2007, QN => n3627);
   KEY_EXPAN0_reg_7_20_inst : FD1 port map( D => n5877, CP => CLK_I, Q => 
                           n_2008, QN => n3614);
   KEY_EXPAN0_reg_6_20_inst : FD1 port map( D => n5876, CP => CLK_I, Q => 
                           n_2009, QN => n3613);
   KEY_EXPAN0_reg_5_20_inst : FD1 port map( D => n5875, CP => CLK_I, Q => 
                           n_2010, QN => n3616);
   KEY_EXPAN0_reg_4_20_inst : FD1 port map( D => n5874, CP => CLK_I, Q => 
                           n_2011, QN => n3615);
   KEY_EXPAN0_reg_3_20_inst : FD1 port map( D => n5873, CP => CLK_I, Q => 
                           n_2012, QN => n3618);
   KEY_EXPAN0_reg_2_20_inst : FD1 port map( D => n5872, CP => CLK_I, Q => 
                           n_2013, QN => n3617);
   KEY_EXPAN0_reg_1_20_inst : FD1 port map( D => n5871, CP => CLK_I, Q => 
                           n_2014, QN => n3620);
   KEY_EXPAN0_reg_0_20_inst : FD1 port map( D => n5870, CP => CLK_I, Q => 
                           n_2015, QN => n3619);
   v_KEY_COL_OUT0_reg_20_inst : FD1 port map( D => n4566, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_20_port, QN => n1906);
   v_TEMP_VECTOR_reg_12_inst : FD1 port map( D => n6683, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_12_port, QN => n_2016);
   KEY_EXPAN0_reg_63_12_inst : FD1 port map( D => n5421, CP => CLK_I, Q => 
                           n_2017, QN => n3542);
   KEY_EXPAN0_reg_62_12_inst : FD1 port map( D => n5420, CP => CLK_I, Q => 
                           n_2018, QN => n3541);
   KEY_EXPAN0_reg_61_12_inst : FD1 port map( D => n5419, CP => CLK_I, Q => 
                           n_2019, QN => n3544);
   KEY_EXPAN0_reg_60_12_inst : FD1 port map( D => n5418, CP => CLK_I, Q => 
                           n_2020, QN => n3543);
   KEY_EXPAN0_reg_59_12_inst : FD1 port map( D => n5417, CP => CLK_I, Q => 
                           n_2021, QN => n3546);
   KEY_EXPAN0_reg_58_12_inst : FD1 port map( D => n5416, CP => CLK_I, Q => 
                           n_2022, QN => n3545);
   KEY_EXPAN0_reg_57_12_inst : FD1 port map( D => n5415, CP => CLK_I, Q => 
                           n_2023, QN => n3548);
   KEY_EXPAN0_reg_56_12_inst : FD1 port map( D => n5414, CP => CLK_I, Q => 
                           n_2024, QN => n3547);
   KEY_EXPAN0_reg_55_12_inst : FD1 port map( D => n5413, CP => CLK_I, Q => 
                           n_2025, QN => n3534);
   KEY_EXPAN0_reg_54_12_inst : FD1 port map( D => n5412, CP => CLK_I, Q => 
                           n_2026, QN => n3533);
   KEY_EXPAN0_reg_53_12_inst : FD1 port map( D => n5411, CP => CLK_I, Q => 
                           n_2027, QN => n3536);
   KEY_EXPAN0_reg_52_12_inst : FD1 port map( D => n5410, CP => CLK_I, Q => 
                           n_2028, QN => n3535);
   KEY_EXPAN0_reg_51_12_inst : FD1 port map( D => n5409, CP => CLK_I, Q => 
                           n_2029, QN => n3538);
   KEY_EXPAN0_reg_50_12_inst : FD1 port map( D => n5408, CP => CLK_I, Q => 
                           n_2030, QN => n3537);
   KEY_EXPAN0_reg_49_12_inst : FD1 port map( D => n5407, CP => CLK_I, Q => 
                           n_2031, QN => n3540);
   KEY_EXPAN0_reg_48_12_inst : FD1 port map( D => n5406, CP => CLK_I, Q => 
                           n_2032, QN => n3539);
   KEY_EXPAN0_reg_47_12_inst : FD1 port map( D => n5405, CP => CLK_I, Q => 
                           n_2033, QN => n3526);
   KEY_EXPAN0_reg_46_12_inst : FD1 port map( D => n5404, CP => CLK_I, Q => 
                           n_2034, QN => n3525);
   KEY_EXPAN0_reg_45_12_inst : FD1 port map( D => n5403, CP => CLK_I, Q => 
                           n_2035, QN => n3528);
   KEY_EXPAN0_reg_44_12_inst : FD1 port map( D => n5402, CP => CLK_I, Q => 
                           n_2036, QN => n3527);
   KEY_EXPAN0_reg_43_12_inst : FD1 port map( D => n5401, CP => CLK_I, Q => 
                           n_2037, QN => n3530);
   KEY_EXPAN0_reg_42_12_inst : FD1 port map( D => n5400, CP => CLK_I, Q => 
                           n_2038, QN => n3529);
   KEY_EXPAN0_reg_41_12_inst : FD1 port map( D => n5399, CP => CLK_I, Q => 
                           n_2039, QN => n3532);
   KEY_EXPAN0_reg_40_12_inst : FD1 port map( D => n5398, CP => CLK_I, Q => 
                           n_2040, QN => n3531);
   KEY_EXPAN0_reg_39_12_inst : FD1 port map( D => n5397, CP => CLK_I, Q => 
                           n_2041, QN => n3518);
   KEY_EXPAN0_reg_38_12_inst : FD1 port map( D => n5396, CP => CLK_I, Q => 
                           n_2042, QN => n3517);
   KEY_EXPAN0_reg_37_12_inst : FD1 port map( D => n5395, CP => CLK_I, Q => 
                           n_2043, QN => n3520);
   KEY_EXPAN0_reg_36_12_inst : FD1 port map( D => n5394, CP => CLK_I, Q => 
                           n_2044, QN => n3519);
   KEY_EXPAN0_reg_35_12_inst : FD1 port map( D => n5393, CP => CLK_I, Q => 
                           n_2045, QN => n3522);
   KEY_EXPAN0_reg_34_12_inst : FD1 port map( D => n5392, CP => CLK_I, Q => 
                           n_2046, QN => n3521);
   KEY_EXPAN0_reg_33_12_inst : FD1 port map( D => n5391, CP => CLK_I, Q => 
                           n_2047, QN => n3524);
   KEY_EXPAN0_reg_32_12_inst : FD1 port map( D => n5390, CP => CLK_I, Q => 
                           n_2048, QN => n3523);
   KEY_EXPAN0_reg_31_12_inst : FD1 port map( D => n5389, CP => CLK_I, Q => 
                           n_2049, QN => n3574);
   KEY_EXPAN0_reg_30_12_inst : FD1 port map( D => n5388, CP => CLK_I, Q => 
                           n_2050, QN => n3573);
   KEY_EXPAN0_reg_29_12_inst : FD1 port map( D => n5387, CP => CLK_I, Q => 
                           n_2051, QN => n3576);
   KEY_EXPAN0_reg_28_12_inst : FD1 port map( D => n5386, CP => CLK_I, Q => 
                           n_2052, QN => n3575);
   KEY_EXPAN0_reg_27_12_inst : FD1 port map( D => n5385, CP => CLK_I, Q => 
                           n_2053, QN => n3578);
   KEY_EXPAN0_reg_26_12_inst : FD1 port map( D => n5384, CP => CLK_I, Q => 
                           n_2054, QN => n3577);
   KEY_EXPAN0_reg_25_12_inst : FD1 port map( D => n5383, CP => CLK_I, Q => 
                           n_2055, QN => n3580);
   KEY_EXPAN0_reg_24_12_inst : FD1 port map( D => n5382, CP => CLK_I, Q => 
                           n_2056, QN => n3579);
   KEY_EXPAN0_reg_23_12_inst : FD1 port map( D => n5381, CP => CLK_I, Q => 
                           n_2057, QN => n3566);
   KEY_EXPAN0_reg_22_12_inst : FD1 port map( D => n5380, CP => CLK_I, Q => 
                           n_2058, QN => n3565);
   KEY_EXPAN0_reg_21_12_inst : FD1 port map( D => n5379, CP => CLK_I, Q => 
                           n_2059, QN => n3568);
   KEY_EXPAN0_reg_20_12_inst : FD1 port map( D => n5378, CP => CLK_I, Q => 
                           n_2060, QN => n3567);
   KEY_EXPAN0_reg_19_12_inst : FD1 port map( D => n5377, CP => CLK_I, Q => 
                           n_2061, QN => n3570);
   KEY_EXPAN0_reg_18_12_inst : FD1 port map( D => n5376, CP => CLK_I, Q => 
                           n_2062, QN => n3569);
   KEY_EXPAN0_reg_17_12_inst : FD1 port map( D => n5375, CP => CLK_I, Q => 
                           n_2063, QN => n3572);
   KEY_EXPAN0_reg_16_12_inst : FD1 port map( D => n5374, CP => CLK_I, Q => 
                           n_2064, QN => n3571);
   KEY_EXPAN0_reg_15_12_inst : FD1 port map( D => n5373, CP => CLK_I, Q => 
                           n_2065, QN => n3558);
   KEY_EXPAN0_reg_14_12_inst : FD1 port map( D => n5372, CP => CLK_I, Q => 
                           n_2066, QN => n3557);
   KEY_EXPAN0_reg_13_12_inst : FD1 port map( D => n5371, CP => CLK_I, Q => 
                           n_2067, QN => n3560);
   KEY_EXPAN0_reg_12_12_inst : FD1 port map( D => n5370, CP => CLK_I, Q => 
                           n_2068, QN => n3559);
   KEY_EXPAN0_reg_11_12_inst : FD1 port map( D => n5369, CP => CLK_I, Q => 
                           n_2069, QN => n3562);
   KEY_EXPAN0_reg_10_12_inst : FD1 port map( D => n5368, CP => CLK_I, Q => 
                           n_2070, QN => n3561);
   KEY_EXPAN0_reg_9_12_inst : FD1 port map( D => n5367, CP => CLK_I, Q => 
                           n_2071, QN => n3564);
   KEY_EXPAN0_reg_8_12_inst : FD1 port map( D => n5366, CP => CLK_I, Q => 
                           n_2072, QN => n3563);
   KEY_EXPAN0_reg_7_12_inst : FD1 port map( D => n5365, CP => CLK_I, Q => 
                           n_2073, QN => n3550);
   KEY_EXPAN0_reg_6_12_inst : FD1 port map( D => n5364, CP => CLK_I, Q => 
                           n_2074, QN => n3549);
   KEY_EXPAN0_reg_5_12_inst : FD1 port map( D => n5363, CP => CLK_I, Q => 
                           n_2075, QN => n3552);
   KEY_EXPAN0_reg_4_12_inst : FD1 port map( D => n5362, CP => CLK_I, Q => 
                           n_2076, QN => n3551);
   KEY_EXPAN0_reg_3_12_inst : FD1 port map( D => n5361, CP => CLK_I, Q => 
                           n_2077, QN => n3554);
   KEY_EXPAN0_reg_2_12_inst : FD1 port map( D => n5360, CP => CLK_I, Q => 
                           n_2078, QN => n3553);
   KEY_EXPAN0_reg_1_12_inst : FD1 port map( D => n5359, CP => CLK_I, Q => 
                           n_2079, QN => n3556);
   KEY_EXPAN0_reg_0_12_inst : FD1 port map( D => n5358, CP => CLK_I, Q => 
                           n_2080, QN => n3555);
   v_KEY_COL_OUT0_reg_12_inst : FD1 port map( D => n4565, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_12_port, QN => n1904);
   v_TEMP_VECTOR_reg_3_inst : FD1 port map( D => n6692, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_3_port, QN => n_2081);
   KEY_EXPAN0_reg_63_3_inst : FD1 port map( D => n4845, CP => CLK_I, Q => 
                           n_2082, QN => n3478);
   KEY_EXPAN0_reg_62_3_inst : FD1 port map( D => n4844, CP => CLK_I, Q => 
                           n_2083, QN => n3477);
   KEY_EXPAN0_reg_61_3_inst : FD1 port map( D => n4843, CP => CLK_I, Q => 
                           n_2084, QN => n3480);
   KEY_EXPAN0_reg_60_3_inst : FD1 port map( D => n4842, CP => CLK_I, Q => 
                           n_2085, QN => n3479);
   KEY_EXPAN0_reg_59_3_inst : FD1 port map( D => n4841, CP => CLK_I, Q => 
                           n_2086, QN => n3482);
   KEY_EXPAN0_reg_58_3_inst : FD1 port map( D => n4840, CP => CLK_I, Q => 
                           n_2087, QN => n3481);
   KEY_EXPAN0_reg_57_3_inst : FD1 port map( D => n4839, CP => CLK_I, Q => 
                           n_2088, QN => n3484);
   KEY_EXPAN0_reg_56_3_inst : FD1 port map( D => n4838, CP => CLK_I, Q => 
                           n_2089, QN => n3483);
   KEY_EXPAN0_reg_55_3_inst : FD1 port map( D => n4837, CP => CLK_I, Q => 
                           n_2090, QN => n3470);
   KEY_EXPAN0_reg_54_3_inst : FD1 port map( D => n4836, CP => CLK_I, Q => 
                           n_2091, QN => n3469);
   KEY_EXPAN0_reg_53_3_inst : FD1 port map( D => n4835, CP => CLK_I, Q => 
                           n_2092, QN => n3472);
   KEY_EXPAN0_reg_52_3_inst : FD1 port map( D => n4834, CP => CLK_I, Q => 
                           n_2093, QN => n3471);
   KEY_EXPAN0_reg_51_3_inst : FD1 port map( D => n4833, CP => CLK_I, Q => 
                           n_2094, QN => n3474);
   KEY_EXPAN0_reg_50_3_inst : FD1 port map( D => n4832, CP => CLK_I, Q => 
                           n_2095, QN => n3473);
   KEY_EXPAN0_reg_49_3_inst : FD1 port map( D => n4831, CP => CLK_I, Q => 
                           n_2096, QN => n3476);
   KEY_EXPAN0_reg_48_3_inst : FD1 port map( D => n4830, CP => CLK_I, Q => 
                           n_2097, QN => n3475);
   KEY_EXPAN0_reg_47_3_inst : FD1 port map( D => n4829, CP => CLK_I, Q => 
                           n_2098, QN => n3462);
   KEY_EXPAN0_reg_46_3_inst : FD1 port map( D => n4828, CP => CLK_I, Q => 
                           n_2099, QN => n3461);
   KEY_EXPAN0_reg_45_3_inst : FD1 port map( D => n4827, CP => CLK_I, Q => 
                           n_2100, QN => n3464);
   KEY_EXPAN0_reg_44_3_inst : FD1 port map( D => n4826, CP => CLK_I, Q => 
                           n_2101, QN => n3463);
   KEY_EXPAN0_reg_43_3_inst : FD1 port map( D => n4825, CP => CLK_I, Q => 
                           n_2102, QN => n3466);
   KEY_EXPAN0_reg_42_3_inst : FD1 port map( D => n4824, CP => CLK_I, Q => 
                           n_2103, QN => n3465);
   KEY_EXPAN0_reg_41_3_inst : FD1 port map( D => n4823, CP => CLK_I, Q => 
                           n_2104, QN => n3468);
   KEY_EXPAN0_reg_40_3_inst : FD1 port map( D => n4822, CP => CLK_I, Q => 
                           n_2105, QN => n3467);
   KEY_EXPAN0_reg_39_3_inst : FD1 port map( D => n4821, CP => CLK_I, Q => 
                           n_2106, QN => n3454);
   KEY_EXPAN0_reg_38_3_inst : FD1 port map( D => n4820, CP => CLK_I, Q => 
                           n_2107, QN => n3453);
   KEY_EXPAN0_reg_37_3_inst : FD1 port map( D => n4819, CP => CLK_I, Q => 
                           n_2108, QN => n3456);
   KEY_EXPAN0_reg_36_3_inst : FD1 port map( D => n4818, CP => CLK_I, Q => 
                           n_2109, QN => n3455);
   KEY_EXPAN0_reg_35_3_inst : FD1 port map( D => n4817, CP => CLK_I, Q => 
                           n_2110, QN => n3458);
   KEY_EXPAN0_reg_34_3_inst : FD1 port map( D => n4816, CP => CLK_I, Q => 
                           n_2111, QN => n3457);
   KEY_EXPAN0_reg_33_3_inst : FD1 port map( D => n4815, CP => CLK_I, Q => 
                           n_2112, QN => n3460);
   KEY_EXPAN0_reg_32_3_inst : FD1 port map( D => n4814, CP => CLK_I, Q => 
                           n_2113, QN => n3459);
   KEY_EXPAN0_reg_31_3_inst : FD1 port map( D => n4813, CP => CLK_I, Q => 
                           n_2114, QN => n3510);
   KEY_EXPAN0_reg_30_3_inst : FD1 port map( D => n4812, CP => CLK_I, Q => 
                           n_2115, QN => n3509);
   KEY_EXPAN0_reg_29_3_inst : FD1 port map( D => n4811, CP => CLK_I, Q => 
                           n_2116, QN => n3512);
   KEY_EXPAN0_reg_28_3_inst : FD1 port map( D => n4810, CP => CLK_I, Q => 
                           n_2117, QN => n3511);
   KEY_EXPAN0_reg_27_3_inst : FD1 port map( D => n4809, CP => CLK_I, Q => 
                           n_2118, QN => n3514);
   KEY_EXPAN0_reg_26_3_inst : FD1 port map( D => n4808, CP => CLK_I, Q => 
                           n_2119, QN => n3513);
   KEY_EXPAN0_reg_25_3_inst : FD1 port map( D => n4807, CP => CLK_I, Q => 
                           n_2120, QN => n3516);
   KEY_EXPAN0_reg_24_3_inst : FD1 port map( D => n4806, CP => CLK_I, Q => 
                           n_2121, QN => n3515);
   KEY_EXPAN0_reg_23_3_inst : FD1 port map( D => n4805, CP => CLK_I, Q => 
                           n_2122, QN => n3502);
   KEY_EXPAN0_reg_22_3_inst : FD1 port map( D => n4804, CP => CLK_I, Q => 
                           n_2123, QN => n3501);
   KEY_EXPAN0_reg_21_3_inst : FD1 port map( D => n4803, CP => CLK_I, Q => 
                           n_2124, QN => n3504);
   KEY_EXPAN0_reg_20_3_inst : FD1 port map( D => n4802, CP => CLK_I, Q => 
                           n_2125, QN => n3503);
   KEY_EXPAN0_reg_19_3_inst : FD1 port map( D => n4801, CP => CLK_I, Q => 
                           n_2126, QN => n3506);
   KEY_EXPAN0_reg_18_3_inst : FD1 port map( D => n4800, CP => CLK_I, Q => 
                           n_2127, QN => n3505);
   KEY_EXPAN0_reg_17_3_inst : FD1 port map( D => n4799, CP => CLK_I, Q => 
                           n_2128, QN => n3508);
   KEY_EXPAN0_reg_16_3_inst : FD1 port map( D => n4798, CP => CLK_I, Q => 
                           n_2129, QN => n3507);
   KEY_EXPAN0_reg_15_3_inst : FD1 port map( D => n4797, CP => CLK_I, Q => 
                           n_2130, QN => n3494);
   KEY_EXPAN0_reg_14_3_inst : FD1 port map( D => n4796, CP => CLK_I, Q => 
                           n_2131, QN => n3493);
   KEY_EXPAN0_reg_13_3_inst : FD1 port map( D => n4795, CP => CLK_I, Q => 
                           n_2132, QN => n3496);
   KEY_EXPAN0_reg_12_3_inst : FD1 port map( D => n4794, CP => CLK_I, Q => 
                           n_2133, QN => n3495);
   KEY_EXPAN0_reg_11_3_inst : FD1 port map( D => n4793, CP => CLK_I, Q => 
                           n_2134, QN => n3498);
   KEY_EXPAN0_reg_10_3_inst : FD1 port map( D => n4792, CP => CLK_I, Q => 
                           n_2135, QN => n3497);
   KEY_EXPAN0_reg_9_3_inst : FD1 port map( D => n4791, CP => CLK_I, Q => n_2136
                           , QN => n3500);
   KEY_EXPAN0_reg_8_3_inst : FD1 port map( D => n4790, CP => CLK_I, Q => n_2137
                           , QN => n3499);
   KEY_EXPAN0_reg_7_3_inst : FD1 port map( D => n4789, CP => CLK_I, Q => n_2138
                           , QN => n3486);
   KEY_EXPAN0_reg_6_3_inst : FD1 port map( D => n4788, CP => CLK_I, Q => n_2139
                           , QN => n3485);
   KEY_EXPAN0_reg_5_3_inst : FD1 port map( D => n4787, CP => CLK_I, Q => n_2140
                           , QN => n3488);
   KEY_EXPAN0_reg_4_3_inst : FD1 port map( D => n4786, CP => CLK_I, Q => n_2141
                           , QN => n3487);
   KEY_EXPAN0_reg_3_3_inst : FD1 port map( D => n4785, CP => CLK_I, Q => n_2142
                           , QN => n3490);
   KEY_EXPAN0_reg_2_3_inst : FD1 port map( D => n4784, CP => CLK_I, Q => n_2143
                           , QN => n3489);
   KEY_EXPAN0_reg_1_3_inst : FD1 port map( D => n4783, CP => CLK_I, Q => n_2144
                           , QN => n3492);
   KEY_EXPAN0_reg_0_3_inst : FD1 port map( D => n4782, CP => CLK_I, Q => n_2145
                           , QN => n3491);
   v_KEY_COL_OUT0_reg_3_inst : FD1 port map( D => n4564, CP => CLK_I, Q => 
                           n_2146, QN => n1586);
   v_TEMP_VECTOR_reg_27_inst : FD1 port map( D => n6668, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_27_port, QN => n_2147);
   KEY_EXPAN0_reg_63_27_inst : FD1 port map( D => n6381, CP => CLK_I, Q => 
                           n_2148, QN => n3414);
   KEY_EXPAN0_reg_62_27_inst : FD1 port map( D => n6380, CP => CLK_I, Q => 
                           n_2149, QN => n3413);
   KEY_EXPAN0_reg_61_27_inst : FD1 port map( D => n6379, CP => CLK_I, Q => 
                           n_2150, QN => n3416);
   KEY_EXPAN0_reg_60_27_inst : FD1 port map( D => n6378, CP => CLK_I, Q => 
                           n_2151, QN => n3415);
   KEY_EXPAN0_reg_59_27_inst : FD1 port map( D => n6377, CP => CLK_I, Q => 
                           n_2152, QN => n3418);
   KEY_EXPAN0_reg_58_27_inst : FD1 port map( D => n6376, CP => CLK_I, Q => 
                           n_2153, QN => n3417);
   KEY_EXPAN0_reg_57_27_inst : FD1 port map( D => n6375, CP => CLK_I, Q => 
                           n_2154, QN => n3420);
   KEY_EXPAN0_reg_56_27_inst : FD1 port map( D => n6374, CP => CLK_I, Q => 
                           n_2155, QN => n3419);
   KEY_EXPAN0_reg_55_27_inst : FD1 port map( D => n6373, CP => CLK_I, Q => 
                           n_2156, QN => n3406);
   KEY_EXPAN0_reg_54_27_inst : FD1 port map( D => n6372, CP => CLK_I, Q => 
                           n_2157, QN => n3405);
   KEY_EXPAN0_reg_53_27_inst : FD1 port map( D => n6371, CP => CLK_I, Q => 
                           n_2158, QN => n3408);
   KEY_EXPAN0_reg_52_27_inst : FD1 port map( D => n6370, CP => CLK_I, Q => 
                           n_2159, QN => n3407);
   KEY_EXPAN0_reg_51_27_inst : FD1 port map( D => n6369, CP => CLK_I, Q => 
                           n_2160, QN => n3410);
   KEY_EXPAN0_reg_50_27_inst : FD1 port map( D => n6368, CP => CLK_I, Q => 
                           n_2161, QN => n3409);
   KEY_EXPAN0_reg_49_27_inst : FD1 port map( D => n6367, CP => CLK_I, Q => 
                           n_2162, QN => n3412);
   KEY_EXPAN0_reg_48_27_inst : FD1 port map( D => n6366, CP => CLK_I, Q => 
                           n_2163, QN => n3411);
   KEY_EXPAN0_reg_47_27_inst : FD1 port map( D => n6365, CP => CLK_I, Q => 
                           n_2164, QN => n3398);
   KEY_EXPAN0_reg_46_27_inst : FD1 port map( D => n6364, CP => CLK_I, Q => 
                           n_2165, QN => n3397);
   KEY_EXPAN0_reg_45_27_inst : FD1 port map( D => n6363, CP => CLK_I, Q => 
                           n_2166, QN => n3400);
   KEY_EXPAN0_reg_44_27_inst : FD1 port map( D => n6362, CP => CLK_I, Q => 
                           n_2167, QN => n3399);
   KEY_EXPAN0_reg_43_27_inst : FD1 port map( D => n6361, CP => CLK_I, Q => 
                           n_2168, QN => n3402);
   KEY_EXPAN0_reg_42_27_inst : FD1 port map( D => n6360, CP => CLK_I, Q => 
                           n_2169, QN => n3401);
   KEY_EXPAN0_reg_41_27_inst : FD1 port map( D => n6359, CP => CLK_I, Q => 
                           n_2170, QN => n3404);
   KEY_EXPAN0_reg_40_27_inst : FD1 port map( D => n6358, CP => CLK_I, Q => 
                           n_2171, QN => n3403);
   KEY_EXPAN0_reg_39_27_inst : FD1 port map( D => n6357, CP => CLK_I, Q => 
                           n_2172, QN => n3390);
   KEY_EXPAN0_reg_38_27_inst : FD1 port map( D => n6356, CP => CLK_I, Q => 
                           n_2173, QN => n3389);
   KEY_EXPAN0_reg_37_27_inst : FD1 port map( D => n6355, CP => CLK_I, Q => 
                           n_2174, QN => n3392);
   KEY_EXPAN0_reg_36_27_inst : FD1 port map( D => n6354, CP => CLK_I, Q => 
                           n_2175, QN => n3391);
   KEY_EXPAN0_reg_35_27_inst : FD1 port map( D => n6353, CP => CLK_I, Q => 
                           n_2176, QN => n3394);
   KEY_EXPAN0_reg_34_27_inst : FD1 port map( D => n6352, CP => CLK_I, Q => 
                           n_2177, QN => n3393);
   KEY_EXPAN0_reg_33_27_inst : FD1 port map( D => n6351, CP => CLK_I, Q => 
                           n_2178, QN => n3396);
   KEY_EXPAN0_reg_32_27_inst : FD1 port map( D => n6350, CP => CLK_I, Q => 
                           n_2179, QN => n3395);
   KEY_EXPAN0_reg_31_27_inst : FD1 port map( D => n6349, CP => CLK_I, Q => 
                           n_2180, QN => n3446);
   KEY_EXPAN0_reg_30_27_inst : FD1 port map( D => n6348, CP => CLK_I, Q => 
                           n_2181, QN => n3445);
   KEY_EXPAN0_reg_29_27_inst : FD1 port map( D => n6347, CP => CLK_I, Q => 
                           n_2182, QN => n3448);
   KEY_EXPAN0_reg_28_27_inst : FD1 port map( D => n6346, CP => CLK_I, Q => 
                           n_2183, QN => n3447);
   KEY_EXPAN0_reg_27_27_inst : FD1 port map( D => n6345, CP => CLK_I, Q => 
                           n_2184, QN => n3450);
   KEY_EXPAN0_reg_26_27_inst : FD1 port map( D => n6344, CP => CLK_I, Q => 
                           n_2185, QN => n3449);
   KEY_EXPAN0_reg_25_27_inst : FD1 port map( D => n6343, CP => CLK_I, Q => 
                           n_2186, QN => n3452);
   KEY_EXPAN0_reg_24_27_inst : FD1 port map( D => n6342, CP => CLK_I, Q => 
                           n_2187, QN => n3451);
   KEY_EXPAN0_reg_23_27_inst : FD1 port map( D => n6341, CP => CLK_I, Q => 
                           n_2188, QN => n3438);
   KEY_EXPAN0_reg_22_27_inst : FD1 port map( D => n6340, CP => CLK_I, Q => 
                           n_2189, QN => n3437);
   KEY_EXPAN0_reg_21_27_inst : FD1 port map( D => n6339, CP => CLK_I, Q => 
                           n_2190, QN => n3440);
   KEY_EXPAN0_reg_20_27_inst : FD1 port map( D => n6338, CP => CLK_I, Q => 
                           n_2191, QN => n3439);
   KEY_EXPAN0_reg_19_27_inst : FD1 port map( D => n6337, CP => CLK_I, Q => 
                           n_2192, QN => n3442);
   KEY_EXPAN0_reg_18_27_inst : FD1 port map( D => n6336, CP => CLK_I, Q => 
                           n_2193, QN => n3441);
   KEY_EXPAN0_reg_17_27_inst : FD1 port map( D => n6335, CP => CLK_I, Q => 
                           n_2194, QN => n3444);
   KEY_EXPAN0_reg_16_27_inst : FD1 port map( D => n6334, CP => CLK_I, Q => 
                           n_2195, QN => n3443);
   KEY_EXPAN0_reg_15_27_inst : FD1 port map( D => n6333, CP => CLK_I, Q => 
                           n_2196, QN => n3430);
   KEY_EXPAN0_reg_14_27_inst : FD1 port map( D => n6332, CP => CLK_I, Q => 
                           n_2197, QN => n3429);
   KEY_EXPAN0_reg_13_27_inst : FD1 port map( D => n6331, CP => CLK_I, Q => 
                           n_2198, QN => n3432);
   KEY_EXPAN0_reg_12_27_inst : FD1 port map( D => n6330, CP => CLK_I, Q => 
                           n_2199, QN => n3431);
   KEY_EXPAN0_reg_11_27_inst : FD1 port map( D => n6329, CP => CLK_I, Q => 
                           n_2200, QN => n3434);
   KEY_EXPAN0_reg_10_27_inst : FD1 port map( D => n6328, CP => CLK_I, Q => 
                           n_2201, QN => n3433);
   KEY_EXPAN0_reg_9_27_inst : FD1 port map( D => n6327, CP => CLK_I, Q => 
                           n_2202, QN => n3436);
   KEY_EXPAN0_reg_8_27_inst : FD1 port map( D => n6326, CP => CLK_I, Q => 
                           n_2203, QN => n3435);
   KEY_EXPAN0_reg_7_27_inst : FD1 port map( D => n6325, CP => CLK_I, Q => 
                           n_2204, QN => n3422);
   KEY_EXPAN0_reg_6_27_inst : FD1 port map( D => n6324, CP => CLK_I, Q => 
                           n_2205, QN => n3421);
   KEY_EXPAN0_reg_5_27_inst : FD1 port map( D => n6323, CP => CLK_I, Q => 
                           n_2206, QN => n3424);
   KEY_EXPAN0_reg_4_27_inst : FD1 port map( D => n6322, CP => CLK_I, Q => 
                           n_2207, QN => n3423);
   KEY_EXPAN0_reg_3_27_inst : FD1 port map( D => n6321, CP => CLK_I, Q => 
                           n_2208, QN => n3426);
   KEY_EXPAN0_reg_2_27_inst : FD1 port map( D => n6320, CP => CLK_I, Q => 
                           n_2209, QN => n3425);
   KEY_EXPAN0_reg_1_27_inst : FD1 port map( D => n6319, CP => CLK_I, Q => 
                           n_2210, QN => n3428);
   KEY_EXPAN0_reg_0_27_inst : FD1 port map( D => n6318, CP => CLK_I, Q => 
                           n_2211, QN => n3427);
   v_KEY_COL_OUT0_reg_27_inst : FD1 port map( D => n4563, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_27_port, QN => n357);
   v_TEMP_VECTOR_reg_19_inst : FD1 port map( D => n6676, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_19_port, QN => n_2212);
   KEY_EXPAN0_reg_63_19_inst : FD1 port map( D => n5869, CP => CLK_I, Q => 
                           n_2213, QN => n3350);
   KEY_EXPAN0_reg_62_19_inst : FD1 port map( D => n5868, CP => CLK_I, Q => 
                           n_2214, QN => n3349);
   KEY_EXPAN0_reg_61_19_inst : FD1 port map( D => n5867, CP => CLK_I, Q => 
                           n_2215, QN => n3352);
   KEY_EXPAN0_reg_60_19_inst : FD1 port map( D => n5866, CP => CLK_I, Q => 
                           n_2216, QN => n3351);
   KEY_EXPAN0_reg_59_19_inst : FD1 port map( D => n5865, CP => CLK_I, Q => 
                           n_2217, QN => n3354);
   KEY_EXPAN0_reg_58_19_inst : FD1 port map( D => n5864, CP => CLK_I, Q => 
                           n_2218, QN => n3353);
   KEY_EXPAN0_reg_57_19_inst : FD1 port map( D => n5863, CP => CLK_I, Q => 
                           n_2219, QN => n3356);
   KEY_EXPAN0_reg_56_19_inst : FD1 port map( D => n5862, CP => CLK_I, Q => 
                           n_2220, QN => n3355);
   KEY_EXPAN0_reg_55_19_inst : FD1 port map( D => n5861, CP => CLK_I, Q => 
                           n_2221, QN => n3342);
   KEY_EXPAN0_reg_54_19_inst : FD1 port map( D => n5860, CP => CLK_I, Q => 
                           n_2222, QN => n3341);
   KEY_EXPAN0_reg_53_19_inst : FD1 port map( D => n5859, CP => CLK_I, Q => 
                           n_2223, QN => n3344);
   KEY_EXPAN0_reg_52_19_inst : FD1 port map( D => n5858, CP => CLK_I, Q => 
                           n_2224, QN => n3343);
   KEY_EXPAN0_reg_51_19_inst : FD1 port map( D => n5857, CP => CLK_I, Q => 
                           n_2225, QN => n3346);
   KEY_EXPAN0_reg_50_19_inst : FD1 port map( D => n5856, CP => CLK_I, Q => 
                           n_2226, QN => n3345);
   KEY_EXPAN0_reg_49_19_inst : FD1 port map( D => n5855, CP => CLK_I, Q => 
                           n_2227, QN => n3348);
   KEY_EXPAN0_reg_48_19_inst : FD1 port map( D => n5854, CP => CLK_I, Q => 
                           n_2228, QN => n3347);
   KEY_EXPAN0_reg_47_19_inst : FD1 port map( D => n5853, CP => CLK_I, Q => 
                           n_2229, QN => n3334);
   KEY_EXPAN0_reg_46_19_inst : FD1 port map( D => n5852, CP => CLK_I, Q => 
                           n_2230, QN => n3333);
   KEY_EXPAN0_reg_45_19_inst : FD1 port map( D => n5851, CP => CLK_I, Q => 
                           n_2231, QN => n3336);
   KEY_EXPAN0_reg_44_19_inst : FD1 port map( D => n5850, CP => CLK_I, Q => 
                           n_2232, QN => n3335);
   KEY_EXPAN0_reg_43_19_inst : FD1 port map( D => n5849, CP => CLK_I, Q => 
                           n_2233, QN => n3338);
   KEY_EXPAN0_reg_42_19_inst : FD1 port map( D => n5848, CP => CLK_I, Q => 
                           n_2234, QN => n3337);
   KEY_EXPAN0_reg_41_19_inst : FD1 port map( D => n5847, CP => CLK_I, Q => 
                           n_2235, QN => n3340);
   KEY_EXPAN0_reg_40_19_inst : FD1 port map( D => n5846, CP => CLK_I, Q => 
                           n_2236, QN => n3339);
   KEY_EXPAN0_reg_39_19_inst : FD1 port map( D => n5845, CP => CLK_I, Q => 
                           n_2237, QN => n3326);
   KEY_EXPAN0_reg_38_19_inst : FD1 port map( D => n5844, CP => CLK_I, Q => 
                           n_2238, QN => n3325);
   KEY_EXPAN0_reg_37_19_inst : FD1 port map( D => n5843, CP => CLK_I, Q => 
                           n_2239, QN => n3328);
   KEY_EXPAN0_reg_36_19_inst : FD1 port map( D => n5842, CP => CLK_I, Q => 
                           n_2240, QN => n3327);
   KEY_EXPAN0_reg_35_19_inst : FD1 port map( D => n5841, CP => CLK_I, Q => 
                           n_2241, QN => n3330);
   KEY_EXPAN0_reg_34_19_inst : FD1 port map( D => n5840, CP => CLK_I, Q => 
                           n_2242, QN => n3329);
   KEY_EXPAN0_reg_33_19_inst : FD1 port map( D => n5839, CP => CLK_I, Q => 
                           n_2243, QN => n3332);
   KEY_EXPAN0_reg_32_19_inst : FD1 port map( D => n5838, CP => CLK_I, Q => 
                           n_2244, QN => n3331);
   KEY_EXPAN0_reg_31_19_inst : FD1 port map( D => n5837, CP => CLK_I, Q => 
                           n_2245, QN => n3382);
   KEY_EXPAN0_reg_30_19_inst : FD1 port map( D => n5836, CP => CLK_I, Q => 
                           n_2246, QN => n3381);
   KEY_EXPAN0_reg_29_19_inst : FD1 port map( D => n5835, CP => CLK_I, Q => 
                           n_2247, QN => n3384);
   KEY_EXPAN0_reg_28_19_inst : FD1 port map( D => n5834, CP => CLK_I, Q => 
                           n_2248, QN => n3383);
   KEY_EXPAN0_reg_27_19_inst : FD1 port map( D => n5833, CP => CLK_I, Q => 
                           n_2249, QN => n3386);
   KEY_EXPAN0_reg_26_19_inst : FD1 port map( D => n5832, CP => CLK_I, Q => 
                           n_2250, QN => n3385);
   KEY_EXPAN0_reg_25_19_inst : FD1 port map( D => n5831, CP => CLK_I, Q => 
                           n_2251, QN => n3388);
   KEY_EXPAN0_reg_24_19_inst : FD1 port map( D => n5830, CP => CLK_I, Q => 
                           n_2252, QN => n3387);
   KEY_EXPAN0_reg_23_19_inst : FD1 port map( D => n5829, CP => CLK_I, Q => 
                           n_2253, QN => n3374);
   KEY_EXPAN0_reg_22_19_inst : FD1 port map( D => n5828, CP => CLK_I, Q => 
                           n_2254, QN => n3373);
   KEY_EXPAN0_reg_21_19_inst : FD1 port map( D => n5827, CP => CLK_I, Q => 
                           n_2255, QN => n3376);
   KEY_EXPAN0_reg_20_19_inst : FD1 port map( D => n5826, CP => CLK_I, Q => 
                           n_2256, QN => n3375);
   KEY_EXPAN0_reg_19_19_inst : FD1 port map( D => n5825, CP => CLK_I, Q => 
                           n_2257, QN => n3378);
   KEY_EXPAN0_reg_18_19_inst : FD1 port map( D => n5824, CP => CLK_I, Q => 
                           n_2258, QN => n3377);
   KEY_EXPAN0_reg_17_19_inst : FD1 port map( D => n5823, CP => CLK_I, Q => 
                           n_2259, QN => n3380);
   KEY_EXPAN0_reg_16_19_inst : FD1 port map( D => n5822, CP => CLK_I, Q => 
                           n_2260, QN => n3379);
   KEY_EXPAN0_reg_15_19_inst : FD1 port map( D => n5821, CP => CLK_I, Q => 
                           n_2261, QN => n3366);
   KEY_EXPAN0_reg_14_19_inst : FD1 port map( D => n5820, CP => CLK_I, Q => 
                           n_2262, QN => n3365);
   KEY_EXPAN0_reg_13_19_inst : FD1 port map( D => n5819, CP => CLK_I, Q => 
                           n_2263, QN => n3368);
   KEY_EXPAN0_reg_12_19_inst : FD1 port map( D => n5818, CP => CLK_I, Q => 
                           n_2264, QN => n3367);
   KEY_EXPAN0_reg_11_19_inst : FD1 port map( D => n5817, CP => CLK_I, Q => 
                           n_2265, QN => n3370);
   KEY_EXPAN0_reg_10_19_inst : FD1 port map( D => n5816, CP => CLK_I, Q => 
                           n_2266, QN => n3369);
   KEY_EXPAN0_reg_9_19_inst : FD1 port map( D => n5815, CP => CLK_I, Q => 
                           n_2267, QN => n3372);
   KEY_EXPAN0_reg_8_19_inst : FD1 port map( D => n5814, CP => CLK_I, Q => 
                           n_2268, QN => n3371);
   KEY_EXPAN0_reg_7_19_inst : FD1 port map( D => n5813, CP => CLK_I, Q => 
                           n_2269, QN => n3358);
   KEY_EXPAN0_reg_6_19_inst : FD1 port map( D => n5812, CP => CLK_I, Q => 
                           n_2270, QN => n3357);
   KEY_EXPAN0_reg_5_19_inst : FD1 port map( D => n5811, CP => CLK_I, Q => 
                           n_2271, QN => n3360);
   KEY_EXPAN0_reg_4_19_inst : FD1 port map( D => n5810, CP => CLK_I, Q => 
                           n_2272, QN => n3359);
   KEY_EXPAN0_reg_3_19_inst : FD1 port map( D => n5809, CP => CLK_I, Q => 
                           n_2273, QN => n3362);
   KEY_EXPAN0_reg_2_19_inst : FD1 port map( D => n5808, CP => CLK_I, Q => 
                           n_2274, QN => n3361);
   KEY_EXPAN0_reg_1_19_inst : FD1 port map( D => n5807, CP => CLK_I, Q => 
                           n_2275, QN => n3364);
   KEY_EXPAN0_reg_0_19_inst : FD1 port map( D => n5806, CP => CLK_I, Q => 
                           n_2276, QN => n3363);
   v_KEY_COL_OUT0_reg_19_inst : FD1 port map( D => n4562, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_19_port, QN => n1367);
   v_TEMP_VECTOR_reg_11_inst : FD1 port map( D => n6684, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_11_port, QN => n_2277);
   KEY_EXPAN0_reg_63_11_inst : FD1 port map( D => n5357, CP => CLK_I, Q => 
                           n_2278, QN => n3286);
   KEY_EXPAN0_reg_62_11_inst : FD1 port map( D => n5356, CP => CLK_I, Q => 
                           n_2279, QN => n3285);
   KEY_EXPAN0_reg_61_11_inst : FD1 port map( D => n5355, CP => CLK_I, Q => 
                           n_2280, QN => n3288);
   KEY_EXPAN0_reg_60_11_inst : FD1 port map( D => n5354, CP => CLK_I, Q => 
                           n_2281, QN => n3287);
   KEY_EXPAN0_reg_59_11_inst : FD1 port map( D => n5353, CP => CLK_I, Q => 
                           n_2282, QN => n3290);
   KEY_EXPAN0_reg_58_11_inst : FD1 port map( D => n5352, CP => CLK_I, Q => 
                           n_2283, QN => n3289);
   KEY_EXPAN0_reg_57_11_inst : FD1 port map( D => n5351, CP => CLK_I, Q => 
                           n_2284, QN => n3292);
   KEY_EXPAN0_reg_56_11_inst : FD1 port map( D => n5350, CP => CLK_I, Q => 
                           n_2285, QN => n3291);
   KEY_EXPAN0_reg_55_11_inst : FD1 port map( D => n5349, CP => CLK_I, Q => 
                           n_2286, QN => n3278);
   KEY_EXPAN0_reg_54_11_inst : FD1 port map( D => n5348, CP => CLK_I, Q => 
                           n_2287, QN => n3277);
   KEY_EXPAN0_reg_53_11_inst : FD1 port map( D => n5347, CP => CLK_I, Q => 
                           n_2288, QN => n3280);
   KEY_EXPAN0_reg_52_11_inst : FD1 port map( D => n5346, CP => CLK_I, Q => 
                           n_2289, QN => n3279);
   KEY_EXPAN0_reg_51_11_inst : FD1 port map( D => n5345, CP => CLK_I, Q => 
                           n_2290, QN => n3282);
   KEY_EXPAN0_reg_50_11_inst : FD1 port map( D => n5344, CP => CLK_I, Q => 
                           n_2291, QN => n3281);
   KEY_EXPAN0_reg_49_11_inst : FD1 port map( D => n5343, CP => CLK_I, Q => 
                           n_2292, QN => n3284);
   KEY_EXPAN0_reg_48_11_inst : FD1 port map( D => n5342, CP => CLK_I, Q => 
                           n_2293, QN => n3283);
   KEY_EXPAN0_reg_47_11_inst : FD1 port map( D => n5341, CP => CLK_I, Q => 
                           n_2294, QN => n3270);
   KEY_EXPAN0_reg_46_11_inst : FD1 port map( D => n5340, CP => CLK_I, Q => 
                           n_2295, QN => n3269);
   KEY_EXPAN0_reg_45_11_inst : FD1 port map( D => n5339, CP => CLK_I, Q => 
                           n_2296, QN => n3272);
   KEY_EXPAN0_reg_44_11_inst : FD1 port map( D => n5338, CP => CLK_I, Q => 
                           n_2297, QN => n3271);
   KEY_EXPAN0_reg_43_11_inst : FD1 port map( D => n5337, CP => CLK_I, Q => 
                           n_2298, QN => n3274);
   KEY_EXPAN0_reg_42_11_inst : FD1 port map( D => n5336, CP => CLK_I, Q => 
                           n_2299, QN => n3273);
   KEY_EXPAN0_reg_41_11_inst : FD1 port map( D => n5335, CP => CLK_I, Q => 
                           n_2300, QN => n3276);
   KEY_EXPAN0_reg_40_11_inst : FD1 port map( D => n5334, CP => CLK_I, Q => 
                           n_2301, QN => n3275);
   KEY_EXPAN0_reg_39_11_inst : FD1 port map( D => n5333, CP => CLK_I, Q => 
                           n_2302, QN => n3262);
   KEY_EXPAN0_reg_38_11_inst : FD1 port map( D => n5332, CP => CLK_I, Q => 
                           n_2303, QN => n3261);
   KEY_EXPAN0_reg_37_11_inst : FD1 port map( D => n5331, CP => CLK_I, Q => 
                           n_2304, QN => n3264);
   KEY_EXPAN0_reg_36_11_inst : FD1 port map( D => n5330, CP => CLK_I, Q => 
                           n_2305, QN => n3263);
   KEY_EXPAN0_reg_35_11_inst : FD1 port map( D => n5329, CP => CLK_I, Q => 
                           n_2306, QN => n3266);
   KEY_EXPAN0_reg_34_11_inst : FD1 port map( D => n5328, CP => CLK_I, Q => 
                           n_2307, QN => n3265);
   KEY_EXPAN0_reg_33_11_inst : FD1 port map( D => n5327, CP => CLK_I, Q => 
                           n_2308, QN => n3268);
   KEY_EXPAN0_reg_32_11_inst : FD1 port map( D => n5326, CP => CLK_I, Q => 
                           n_2309, QN => n3267);
   KEY_EXPAN0_reg_31_11_inst : FD1 port map( D => n5325, CP => CLK_I, Q => 
                           n_2310, QN => n3318);
   KEY_EXPAN0_reg_30_11_inst : FD1 port map( D => n5324, CP => CLK_I, Q => 
                           n_2311, QN => n3317);
   KEY_EXPAN0_reg_29_11_inst : FD1 port map( D => n5323, CP => CLK_I, Q => 
                           n_2312, QN => n3320);
   KEY_EXPAN0_reg_28_11_inst : FD1 port map( D => n5322, CP => CLK_I, Q => 
                           n_2313, QN => n3319);
   KEY_EXPAN0_reg_27_11_inst : FD1 port map( D => n5321, CP => CLK_I, Q => 
                           n_2314, QN => n3322);
   KEY_EXPAN0_reg_26_11_inst : FD1 port map( D => n5320, CP => CLK_I, Q => 
                           n_2315, QN => n3321);
   KEY_EXPAN0_reg_25_11_inst : FD1 port map( D => n5319, CP => CLK_I, Q => 
                           n_2316, QN => n3324);
   KEY_EXPAN0_reg_24_11_inst : FD1 port map( D => n5318, CP => CLK_I, Q => 
                           n_2317, QN => n3323);
   KEY_EXPAN0_reg_23_11_inst : FD1 port map( D => n5317, CP => CLK_I, Q => 
                           n_2318, QN => n3310);
   KEY_EXPAN0_reg_22_11_inst : FD1 port map( D => n5316, CP => CLK_I, Q => 
                           n_2319, QN => n3309);
   KEY_EXPAN0_reg_21_11_inst : FD1 port map( D => n5315, CP => CLK_I, Q => 
                           n_2320, QN => n3312);
   KEY_EXPAN0_reg_20_11_inst : FD1 port map( D => n5314, CP => CLK_I, Q => 
                           n_2321, QN => n3311);
   KEY_EXPAN0_reg_19_11_inst : FD1 port map( D => n5313, CP => CLK_I, Q => 
                           n_2322, QN => n3314);
   KEY_EXPAN0_reg_18_11_inst : FD1 port map( D => n5312, CP => CLK_I, Q => 
                           n_2323, QN => n3313);
   KEY_EXPAN0_reg_17_11_inst : FD1 port map( D => n5311, CP => CLK_I, Q => 
                           n_2324, QN => n3316);
   KEY_EXPAN0_reg_16_11_inst : FD1 port map( D => n5310, CP => CLK_I, Q => 
                           n_2325, QN => n3315);
   KEY_EXPAN0_reg_15_11_inst : FD1 port map( D => n5309, CP => CLK_I, Q => 
                           n_2326, QN => n3302);
   KEY_EXPAN0_reg_14_11_inst : FD1 port map( D => n5308, CP => CLK_I, Q => 
                           n_2327, QN => n3301);
   KEY_EXPAN0_reg_13_11_inst : FD1 port map( D => n5307, CP => CLK_I, Q => 
                           n_2328, QN => n3304);
   KEY_EXPAN0_reg_12_11_inst : FD1 port map( D => n5306, CP => CLK_I, Q => 
                           n_2329, QN => n3303);
   KEY_EXPAN0_reg_11_11_inst : FD1 port map( D => n5305, CP => CLK_I, Q => 
                           n_2330, QN => n3306);
   KEY_EXPAN0_reg_10_11_inst : FD1 port map( D => n5304, CP => CLK_I, Q => 
                           n_2331, QN => n3305);
   KEY_EXPAN0_reg_9_11_inst : FD1 port map( D => n5303, CP => CLK_I, Q => 
                           n_2332, QN => n3308);
   KEY_EXPAN0_reg_8_11_inst : FD1 port map( D => n5302, CP => CLK_I, Q => 
                           n_2333, QN => n3307);
   KEY_EXPAN0_reg_7_11_inst : FD1 port map( D => n5301, CP => CLK_I, Q => 
                           n_2334, QN => n3294);
   KEY_EXPAN0_reg_6_11_inst : FD1 port map( D => n5300, CP => CLK_I, Q => 
                           n_2335, QN => n3293);
   KEY_EXPAN0_reg_5_11_inst : FD1 port map( D => n5299, CP => CLK_I, Q => 
                           n_2336, QN => n3296);
   KEY_EXPAN0_reg_4_11_inst : FD1 port map( D => n5298, CP => CLK_I, Q => 
                           n_2337, QN => n3295);
   KEY_EXPAN0_reg_3_11_inst : FD1 port map( D => n5297, CP => CLK_I, Q => 
                           n_2338, QN => n3298);
   KEY_EXPAN0_reg_2_11_inst : FD1 port map( D => n5296, CP => CLK_I, Q => 
                           n_2339, QN => n3297);
   KEY_EXPAN0_reg_1_11_inst : FD1 port map( D => n5295, CP => CLK_I, Q => 
                           n_2340, QN => n3300);
   KEY_EXPAN0_reg_0_11_inst : FD1 port map( D => n5294, CP => CLK_I, Q => 
                           n_2341, QN => n3299);
   v_KEY_COL_OUT0_reg_11_inst : FD1 port map( D => n4561, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_11_port, QN => n356);
   v_TEMP_VECTOR_reg_2_inst : FD1 port map( D => n6693, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_2_port, QN => n_2342);
   KEY_EXPAN0_reg_63_2_inst : FD1 port map( D => n4781, CP => CLK_I, Q => 
                           n_2343, QN => n3222);
   KEY_EXPAN0_reg_62_2_inst : FD1 port map( D => n4780, CP => CLK_I, Q => 
                           n_2344, QN => n3221);
   KEY_EXPAN0_reg_61_2_inst : FD1 port map( D => n4779, CP => CLK_I, Q => 
                           n_2345, QN => n3224);
   KEY_EXPAN0_reg_60_2_inst : FD1 port map( D => n4778, CP => CLK_I, Q => 
                           n_2346, QN => n3223);
   KEY_EXPAN0_reg_59_2_inst : FD1 port map( D => n4777, CP => CLK_I, Q => 
                           n_2347, QN => n3226);
   KEY_EXPAN0_reg_58_2_inst : FD1 port map( D => n4776, CP => CLK_I, Q => 
                           n_2348, QN => n3225);
   KEY_EXPAN0_reg_57_2_inst : FD1 port map( D => n4775, CP => CLK_I, Q => 
                           n_2349, QN => n3228);
   KEY_EXPAN0_reg_56_2_inst : FD1 port map( D => n4774, CP => CLK_I, Q => 
                           n_2350, QN => n3227);
   KEY_EXPAN0_reg_55_2_inst : FD1 port map( D => n4773, CP => CLK_I, Q => 
                           n_2351, QN => n3214);
   KEY_EXPAN0_reg_54_2_inst : FD1 port map( D => n4772, CP => CLK_I, Q => 
                           n_2352, QN => n3213);
   KEY_EXPAN0_reg_53_2_inst : FD1 port map( D => n4771, CP => CLK_I, Q => 
                           n_2353, QN => n3216);
   KEY_EXPAN0_reg_52_2_inst : FD1 port map( D => n4770, CP => CLK_I, Q => 
                           n_2354, QN => n3215);
   KEY_EXPAN0_reg_51_2_inst : FD1 port map( D => n4769, CP => CLK_I, Q => 
                           n_2355, QN => n3218);
   KEY_EXPAN0_reg_50_2_inst : FD1 port map( D => n4768, CP => CLK_I, Q => 
                           n_2356, QN => n3217);
   KEY_EXPAN0_reg_49_2_inst : FD1 port map( D => n4767, CP => CLK_I, Q => 
                           n_2357, QN => n3220);
   KEY_EXPAN0_reg_48_2_inst : FD1 port map( D => n4766, CP => CLK_I, Q => 
                           n_2358, QN => n3219);
   KEY_EXPAN0_reg_47_2_inst : FD1 port map( D => n4765, CP => CLK_I, Q => 
                           n_2359, QN => n3206);
   KEY_EXPAN0_reg_46_2_inst : FD1 port map( D => n4764, CP => CLK_I, Q => 
                           n_2360, QN => n3205);
   KEY_EXPAN0_reg_45_2_inst : FD1 port map( D => n4763, CP => CLK_I, Q => 
                           n_2361, QN => n3208);
   KEY_EXPAN0_reg_44_2_inst : FD1 port map( D => n4762, CP => CLK_I, Q => 
                           n_2362, QN => n3207);
   KEY_EXPAN0_reg_43_2_inst : FD1 port map( D => n4761, CP => CLK_I, Q => 
                           n_2363, QN => n3210);
   KEY_EXPAN0_reg_42_2_inst : FD1 port map( D => n4760, CP => CLK_I, Q => 
                           n_2364, QN => n3209);
   KEY_EXPAN0_reg_41_2_inst : FD1 port map( D => n4759, CP => CLK_I, Q => 
                           n_2365, QN => n3212);
   KEY_EXPAN0_reg_40_2_inst : FD1 port map( D => n4758, CP => CLK_I, Q => 
                           n_2366, QN => n3211);
   KEY_EXPAN0_reg_39_2_inst : FD1 port map( D => n4757, CP => CLK_I, Q => 
                           n_2367, QN => n3198);
   KEY_EXPAN0_reg_38_2_inst : FD1 port map( D => n4756, CP => CLK_I, Q => 
                           n_2368, QN => n3197);
   KEY_EXPAN0_reg_37_2_inst : FD1 port map( D => n4755, CP => CLK_I, Q => 
                           n_2369, QN => n3200);
   KEY_EXPAN0_reg_36_2_inst : FD1 port map( D => n4754, CP => CLK_I, Q => 
                           n_2370, QN => n3199);
   KEY_EXPAN0_reg_35_2_inst : FD1 port map( D => n4753, CP => CLK_I, Q => 
                           n_2371, QN => n3202);
   KEY_EXPAN0_reg_34_2_inst : FD1 port map( D => n4752, CP => CLK_I, Q => 
                           n_2372, QN => n3201);
   KEY_EXPAN0_reg_33_2_inst : FD1 port map( D => n4751, CP => CLK_I, Q => 
                           n_2373, QN => n3204);
   KEY_EXPAN0_reg_32_2_inst : FD1 port map( D => n4750, CP => CLK_I, Q => 
                           n_2374, QN => n3203);
   KEY_EXPAN0_reg_31_2_inst : FD1 port map( D => n4749, CP => CLK_I, Q => 
                           n_2375, QN => n3254);
   KEY_EXPAN0_reg_30_2_inst : FD1 port map( D => n4748, CP => CLK_I, Q => 
                           n_2376, QN => n3253);
   KEY_EXPAN0_reg_29_2_inst : FD1 port map( D => n4747, CP => CLK_I, Q => 
                           n_2377, QN => n3256);
   KEY_EXPAN0_reg_28_2_inst : FD1 port map( D => n4746, CP => CLK_I, Q => 
                           n_2378, QN => n3255);
   KEY_EXPAN0_reg_27_2_inst : FD1 port map( D => n4745, CP => CLK_I, Q => 
                           n_2379, QN => n3258);
   KEY_EXPAN0_reg_26_2_inst : FD1 port map( D => n4744, CP => CLK_I, Q => 
                           n_2380, QN => n3257);
   KEY_EXPAN0_reg_25_2_inst : FD1 port map( D => n4743, CP => CLK_I, Q => 
                           n_2381, QN => n3260);
   KEY_EXPAN0_reg_24_2_inst : FD1 port map( D => n4742, CP => CLK_I, Q => 
                           n_2382, QN => n3259);
   KEY_EXPAN0_reg_23_2_inst : FD1 port map( D => n4741, CP => CLK_I, Q => 
                           n_2383, QN => n3246);
   KEY_EXPAN0_reg_22_2_inst : FD1 port map( D => n4740, CP => CLK_I, Q => 
                           n_2384, QN => n3245);
   KEY_EXPAN0_reg_21_2_inst : FD1 port map( D => n4739, CP => CLK_I, Q => 
                           n_2385, QN => n3248);
   KEY_EXPAN0_reg_20_2_inst : FD1 port map( D => n4738, CP => CLK_I, Q => 
                           n_2386, QN => n3247);
   KEY_EXPAN0_reg_19_2_inst : FD1 port map( D => n4737, CP => CLK_I, Q => 
                           n_2387, QN => n3250);
   KEY_EXPAN0_reg_18_2_inst : FD1 port map( D => n4736, CP => CLK_I, Q => 
                           n_2388, QN => n3249);
   KEY_EXPAN0_reg_17_2_inst : FD1 port map( D => n4735, CP => CLK_I, Q => 
                           n_2389, QN => n3252);
   KEY_EXPAN0_reg_16_2_inst : FD1 port map( D => n4734, CP => CLK_I, Q => 
                           n_2390, QN => n3251);
   KEY_EXPAN0_reg_15_2_inst : FD1 port map( D => n4733, CP => CLK_I, Q => 
                           n_2391, QN => n3238);
   KEY_EXPAN0_reg_14_2_inst : FD1 port map( D => n4732, CP => CLK_I, Q => 
                           n_2392, QN => n3237);
   KEY_EXPAN0_reg_13_2_inst : FD1 port map( D => n4731, CP => CLK_I, Q => 
                           n_2393, QN => n3240);
   KEY_EXPAN0_reg_12_2_inst : FD1 port map( D => n4730, CP => CLK_I, Q => 
                           n_2394, QN => n3239);
   KEY_EXPAN0_reg_11_2_inst : FD1 port map( D => n4729, CP => CLK_I, Q => 
                           n_2395, QN => n3242);
   KEY_EXPAN0_reg_10_2_inst : FD1 port map( D => n4728, CP => CLK_I, Q => 
                           n_2396, QN => n3241);
   KEY_EXPAN0_reg_9_2_inst : FD1 port map( D => n4727, CP => CLK_I, Q => n_2397
                           , QN => n3244);
   KEY_EXPAN0_reg_8_2_inst : FD1 port map( D => n4726, CP => CLK_I, Q => n_2398
                           , QN => n3243);
   KEY_EXPAN0_reg_7_2_inst : FD1 port map( D => n4725, CP => CLK_I, Q => n_2399
                           , QN => n3230);
   KEY_EXPAN0_reg_6_2_inst : FD1 port map( D => n4724, CP => CLK_I, Q => n_2400
                           , QN => n3229);
   KEY_EXPAN0_reg_5_2_inst : FD1 port map( D => n4723, CP => CLK_I, Q => n_2401
                           , QN => n3232);
   KEY_EXPAN0_reg_4_2_inst : FD1 port map( D => n4722, CP => CLK_I, Q => n_2402
                           , QN => n3231);
   KEY_EXPAN0_reg_3_2_inst : FD1 port map( D => n4721, CP => CLK_I, Q => n_2403
                           , QN => n3234);
   KEY_EXPAN0_reg_2_2_inst : FD1 port map( D => n4720, CP => CLK_I, Q => n_2404
                           , QN => n3233);
   KEY_EXPAN0_reg_1_2_inst : FD1 port map( D => n4719, CP => CLK_I, Q => n_2405
                           , QN => n3236);
   KEY_EXPAN0_reg_0_2_inst : FD1 port map( D => n4718, CP => CLK_I, Q => n_2406
                           , QN => n3235);
   v_KEY_COL_OUT0_reg_2_inst : FD1 port map( D => n4560, CP => CLK_I, Q => 
                           n_2407, QN => n403);
   v_TEMP_VECTOR_reg_26_inst : FD1 port map( D => n6669, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_26_port, QN => n_2408);
   KEY_EXPAN0_reg_63_26_inst : FD1 port map( D => n6317, CP => CLK_I, Q => 
                           n_2409, QN => n3158);
   KEY_EXPAN0_reg_62_26_inst : FD1 port map( D => n6316, CP => CLK_I, Q => 
                           n_2410, QN => n3157);
   KEY_EXPAN0_reg_61_26_inst : FD1 port map( D => n6315, CP => CLK_I, Q => 
                           n_2411, QN => n3160);
   KEY_EXPAN0_reg_60_26_inst : FD1 port map( D => n6314, CP => CLK_I, Q => 
                           n_2412, QN => n3159);
   KEY_EXPAN0_reg_59_26_inst : FD1 port map( D => n6313, CP => CLK_I, Q => 
                           n_2413, QN => n3162);
   KEY_EXPAN0_reg_58_26_inst : FD1 port map( D => n6312, CP => CLK_I, Q => 
                           n_2414, QN => n3161);
   KEY_EXPAN0_reg_57_26_inst : FD1 port map( D => n6311, CP => CLK_I, Q => 
                           n_2415, QN => n3164);
   KEY_EXPAN0_reg_56_26_inst : FD1 port map( D => n6310, CP => CLK_I, Q => 
                           n_2416, QN => n3163);
   KEY_EXPAN0_reg_55_26_inst : FD1 port map( D => n6309, CP => CLK_I, Q => 
                           n_2417, QN => n3150);
   KEY_EXPAN0_reg_54_26_inst : FD1 port map( D => n6308, CP => CLK_I, Q => 
                           n_2418, QN => n3149);
   KEY_EXPAN0_reg_53_26_inst : FD1 port map( D => n6307, CP => CLK_I, Q => 
                           n_2419, QN => n3152);
   KEY_EXPAN0_reg_52_26_inst : FD1 port map( D => n6306, CP => CLK_I, Q => 
                           n_2420, QN => n3151);
   KEY_EXPAN0_reg_51_26_inst : FD1 port map( D => n6305, CP => CLK_I, Q => 
                           n_2421, QN => n3154);
   KEY_EXPAN0_reg_50_26_inst : FD1 port map( D => n6304, CP => CLK_I, Q => 
                           n_2422, QN => n3153);
   KEY_EXPAN0_reg_49_26_inst : FD1 port map( D => n6303, CP => CLK_I, Q => 
                           n_2423, QN => n3156);
   KEY_EXPAN0_reg_48_26_inst : FD1 port map( D => n6302, CP => CLK_I, Q => 
                           n_2424, QN => n3155);
   KEY_EXPAN0_reg_47_26_inst : FD1 port map( D => n6301, CP => CLK_I, Q => 
                           n_2425, QN => n3142);
   KEY_EXPAN0_reg_46_26_inst : FD1 port map( D => n6300, CP => CLK_I, Q => 
                           n_2426, QN => n3141);
   KEY_EXPAN0_reg_45_26_inst : FD1 port map( D => n6299, CP => CLK_I, Q => 
                           n_2427, QN => n3144);
   KEY_EXPAN0_reg_44_26_inst : FD1 port map( D => n6298, CP => CLK_I, Q => 
                           n_2428, QN => n3143);
   KEY_EXPAN0_reg_43_26_inst : FD1 port map( D => n6297, CP => CLK_I, Q => 
                           n_2429, QN => n3146);
   KEY_EXPAN0_reg_42_26_inst : FD1 port map( D => n6296, CP => CLK_I, Q => 
                           n_2430, QN => n3145);
   KEY_EXPAN0_reg_41_26_inst : FD1 port map( D => n6295, CP => CLK_I, Q => 
                           n_2431, QN => n3148);
   KEY_EXPAN0_reg_40_26_inst : FD1 port map( D => n6294, CP => CLK_I, Q => 
                           n_2432, QN => n3147);
   KEY_EXPAN0_reg_39_26_inst : FD1 port map( D => n6293, CP => CLK_I, Q => 
                           n_2433, QN => n3134);
   KEY_EXPAN0_reg_38_26_inst : FD1 port map( D => n6292, CP => CLK_I, Q => 
                           n_2434, QN => n3133);
   KEY_EXPAN0_reg_37_26_inst : FD1 port map( D => n6291, CP => CLK_I, Q => 
                           n_2435, QN => n3136);
   KEY_EXPAN0_reg_36_26_inst : FD1 port map( D => n6290, CP => CLK_I, Q => 
                           n_2436, QN => n3135);
   KEY_EXPAN0_reg_35_26_inst : FD1 port map( D => n6289, CP => CLK_I, Q => 
                           n_2437, QN => n3138);
   KEY_EXPAN0_reg_34_26_inst : FD1 port map( D => n6288, CP => CLK_I, Q => 
                           n_2438, QN => n3137);
   KEY_EXPAN0_reg_33_26_inst : FD1 port map( D => n6287, CP => CLK_I, Q => 
                           n_2439, QN => n3140);
   KEY_EXPAN0_reg_32_26_inst : FD1 port map( D => n6286, CP => CLK_I, Q => 
                           n_2440, QN => n3139);
   KEY_EXPAN0_reg_31_26_inst : FD1 port map( D => n6285, CP => CLK_I, Q => 
                           n_2441, QN => n3190);
   KEY_EXPAN0_reg_30_26_inst : FD1 port map( D => n6284, CP => CLK_I, Q => 
                           n_2442, QN => n3189);
   KEY_EXPAN0_reg_29_26_inst : FD1 port map( D => n6283, CP => CLK_I, Q => 
                           n_2443, QN => n3192);
   KEY_EXPAN0_reg_28_26_inst : FD1 port map( D => n6282, CP => CLK_I, Q => 
                           n_2444, QN => n3191);
   KEY_EXPAN0_reg_27_26_inst : FD1 port map( D => n6281, CP => CLK_I, Q => 
                           n_2445, QN => n3194);
   KEY_EXPAN0_reg_26_26_inst : FD1 port map( D => n6280, CP => CLK_I, Q => 
                           n_2446, QN => n3193);
   KEY_EXPAN0_reg_25_26_inst : FD1 port map( D => n6279, CP => CLK_I, Q => 
                           n_2447, QN => n3196);
   KEY_EXPAN0_reg_24_26_inst : FD1 port map( D => n6278, CP => CLK_I, Q => 
                           n_2448, QN => n3195);
   KEY_EXPAN0_reg_23_26_inst : FD1 port map( D => n6277, CP => CLK_I, Q => 
                           n_2449, QN => n3182);
   KEY_EXPAN0_reg_22_26_inst : FD1 port map( D => n6276, CP => CLK_I, Q => 
                           n_2450, QN => n3181);
   KEY_EXPAN0_reg_21_26_inst : FD1 port map( D => n6275, CP => CLK_I, Q => 
                           n_2451, QN => n3184);
   KEY_EXPAN0_reg_20_26_inst : FD1 port map( D => n6274, CP => CLK_I, Q => 
                           n_2452, QN => n3183);
   KEY_EXPAN0_reg_19_26_inst : FD1 port map( D => n6273, CP => CLK_I, Q => 
                           n_2453, QN => n3186);
   KEY_EXPAN0_reg_18_26_inst : FD1 port map( D => n6272, CP => CLK_I, Q => 
                           n_2454, QN => n3185);
   KEY_EXPAN0_reg_17_26_inst : FD1 port map( D => n6271, CP => CLK_I, Q => 
                           n_2455, QN => n3188);
   KEY_EXPAN0_reg_16_26_inst : FD1 port map( D => n6270, CP => CLK_I, Q => 
                           n_2456, QN => n3187);
   KEY_EXPAN0_reg_15_26_inst : FD1 port map( D => n6269, CP => CLK_I, Q => 
                           n_2457, QN => n3174);
   KEY_EXPAN0_reg_14_26_inst : FD1 port map( D => n6268, CP => CLK_I, Q => 
                           n_2458, QN => n3173);
   KEY_EXPAN0_reg_13_26_inst : FD1 port map( D => n6267, CP => CLK_I, Q => 
                           n_2459, QN => n3176);
   KEY_EXPAN0_reg_12_26_inst : FD1 port map( D => n6266, CP => CLK_I, Q => 
                           n_2460, QN => n3175);
   KEY_EXPAN0_reg_11_26_inst : FD1 port map( D => n6265, CP => CLK_I, Q => 
                           n_2461, QN => n3178);
   KEY_EXPAN0_reg_10_26_inst : FD1 port map( D => n6264, CP => CLK_I, Q => 
                           n_2462, QN => n3177);
   KEY_EXPAN0_reg_9_26_inst : FD1 port map( D => n6263, CP => CLK_I, Q => 
                           n_2463, QN => n3180);
   KEY_EXPAN0_reg_8_26_inst : FD1 port map( D => n6262, CP => CLK_I, Q => 
                           n_2464, QN => n3179);
   KEY_EXPAN0_reg_7_26_inst : FD1 port map( D => n6261, CP => CLK_I, Q => 
                           n_2465, QN => n3166);
   KEY_EXPAN0_reg_6_26_inst : FD1 port map( D => n6260, CP => CLK_I, Q => 
                           n_2466, QN => n3165);
   KEY_EXPAN0_reg_5_26_inst : FD1 port map( D => n6259, CP => CLK_I, Q => 
                           n_2467, QN => n3168);
   KEY_EXPAN0_reg_4_26_inst : FD1 port map( D => n6258, CP => CLK_I, Q => 
                           n_2468, QN => n3167);
   KEY_EXPAN0_reg_3_26_inst : FD1 port map( D => n6257, CP => CLK_I, Q => 
                           n_2469, QN => n3170);
   KEY_EXPAN0_reg_2_26_inst : FD1 port map( D => n6256, CP => CLK_I, Q => 
                           n_2470, QN => n3169);
   KEY_EXPAN0_reg_1_26_inst : FD1 port map( D => n6255, CP => CLK_I, Q => 
                           n_2471, QN => n3172);
   KEY_EXPAN0_reg_0_26_inst : FD1 port map( D => n6254, CP => CLK_I, Q => 
                           n_2472, QN => n3171);
   v_KEY_COL_OUT0_reg_26_inst : FD1 port map( D => n4559, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_26_port, QN => n391);
   v_TEMP_VECTOR_reg_18_inst : FD1 port map( D => n6677, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_18_port, QN => n_2473);
   KEY_EXPAN0_reg_63_18_inst : FD1 port map( D => n5805, CP => CLK_I, Q => 
                           n_2474, QN => n3094);
   KEY_EXPAN0_reg_62_18_inst : FD1 port map( D => n5804, CP => CLK_I, Q => 
                           n_2475, QN => n3093);
   KEY_EXPAN0_reg_61_18_inst : FD1 port map( D => n5803, CP => CLK_I, Q => 
                           n_2476, QN => n3096);
   KEY_EXPAN0_reg_60_18_inst : FD1 port map( D => n5802, CP => CLK_I, Q => 
                           n_2477, QN => n3095);
   KEY_EXPAN0_reg_59_18_inst : FD1 port map( D => n5801, CP => CLK_I, Q => 
                           n_2478, QN => n3098);
   KEY_EXPAN0_reg_58_18_inst : FD1 port map( D => n5800, CP => CLK_I, Q => 
                           n_2479, QN => n3097);
   KEY_EXPAN0_reg_57_18_inst : FD1 port map( D => n5799, CP => CLK_I, Q => 
                           n_2480, QN => n3100);
   KEY_EXPAN0_reg_56_18_inst : FD1 port map( D => n5798, CP => CLK_I, Q => 
                           n_2481, QN => n3099);
   KEY_EXPAN0_reg_55_18_inst : FD1 port map( D => n5797, CP => CLK_I, Q => 
                           n_2482, QN => n3086);
   KEY_EXPAN0_reg_54_18_inst : FD1 port map( D => n5796, CP => CLK_I, Q => 
                           n_2483, QN => n3085);
   KEY_EXPAN0_reg_53_18_inst : FD1 port map( D => n5795, CP => CLK_I, Q => 
                           n_2484, QN => n3088);
   KEY_EXPAN0_reg_52_18_inst : FD1 port map( D => n5794, CP => CLK_I, Q => 
                           n_2485, QN => n3087);
   KEY_EXPAN0_reg_51_18_inst : FD1 port map( D => n5793, CP => CLK_I, Q => 
                           n_2486, QN => n3090);
   KEY_EXPAN0_reg_50_18_inst : FD1 port map( D => n5792, CP => CLK_I, Q => 
                           n_2487, QN => n3089);
   KEY_EXPAN0_reg_49_18_inst : FD1 port map( D => n5791, CP => CLK_I, Q => 
                           n_2488, QN => n3092);
   KEY_EXPAN0_reg_48_18_inst : FD1 port map( D => n5790, CP => CLK_I, Q => 
                           n_2489, QN => n3091);
   KEY_EXPAN0_reg_47_18_inst : FD1 port map( D => n5789, CP => CLK_I, Q => 
                           n_2490, QN => n3078);
   KEY_EXPAN0_reg_46_18_inst : FD1 port map( D => n5788, CP => CLK_I, Q => 
                           n_2491, QN => n3077);
   KEY_EXPAN0_reg_45_18_inst : FD1 port map( D => n5787, CP => CLK_I, Q => 
                           n_2492, QN => n3080);
   KEY_EXPAN0_reg_44_18_inst : FD1 port map( D => n5786, CP => CLK_I, Q => 
                           n_2493, QN => n3079);
   KEY_EXPAN0_reg_43_18_inst : FD1 port map( D => n5785, CP => CLK_I, Q => 
                           n_2494, QN => n3082);
   KEY_EXPAN0_reg_42_18_inst : FD1 port map( D => n5784, CP => CLK_I, Q => 
                           n_2495, QN => n3081);
   KEY_EXPAN0_reg_41_18_inst : FD1 port map( D => n5783, CP => CLK_I, Q => 
                           n_2496, QN => n3084);
   KEY_EXPAN0_reg_40_18_inst : FD1 port map( D => n5782, CP => CLK_I, Q => 
                           n_2497, QN => n3083);
   KEY_EXPAN0_reg_39_18_inst : FD1 port map( D => n5781, CP => CLK_I, Q => 
                           n_2498, QN => n3070);
   KEY_EXPAN0_reg_38_18_inst : FD1 port map( D => n5780, CP => CLK_I, Q => 
                           n_2499, QN => n3069);
   KEY_EXPAN0_reg_37_18_inst : FD1 port map( D => n5779, CP => CLK_I, Q => 
                           n_2500, QN => n3072);
   KEY_EXPAN0_reg_36_18_inst : FD1 port map( D => n5778, CP => CLK_I, Q => 
                           n_2501, QN => n3071);
   KEY_EXPAN0_reg_35_18_inst : FD1 port map( D => n5777, CP => CLK_I, Q => 
                           n_2502, QN => n3074);
   KEY_EXPAN0_reg_34_18_inst : FD1 port map( D => n5776, CP => CLK_I, Q => 
                           n_2503, QN => n3073);
   KEY_EXPAN0_reg_33_18_inst : FD1 port map( D => n5775, CP => CLK_I, Q => 
                           n_2504, QN => n3076);
   KEY_EXPAN0_reg_32_18_inst : FD1 port map( D => n5774, CP => CLK_I, Q => 
                           n_2505, QN => n3075);
   KEY_EXPAN0_reg_31_18_inst : FD1 port map( D => n5773, CP => CLK_I, Q => 
                           n_2506, QN => n3126);
   KEY_EXPAN0_reg_30_18_inst : FD1 port map( D => n5772, CP => CLK_I, Q => 
                           n_2507, QN => n3125);
   KEY_EXPAN0_reg_29_18_inst : FD1 port map( D => n5771, CP => CLK_I, Q => 
                           n_2508, QN => n3128);
   KEY_EXPAN0_reg_28_18_inst : FD1 port map( D => n5770, CP => CLK_I, Q => 
                           n_2509, QN => n3127);
   KEY_EXPAN0_reg_27_18_inst : FD1 port map( D => n5769, CP => CLK_I, Q => 
                           n_2510, QN => n3130);
   KEY_EXPAN0_reg_26_18_inst : FD1 port map( D => n5768, CP => CLK_I, Q => 
                           n_2511, QN => n3129);
   KEY_EXPAN0_reg_25_18_inst : FD1 port map( D => n5767, CP => CLK_I, Q => 
                           n_2512, QN => n3132);
   KEY_EXPAN0_reg_24_18_inst : FD1 port map( D => n5766, CP => CLK_I, Q => 
                           n_2513, QN => n3131);
   KEY_EXPAN0_reg_23_18_inst : FD1 port map( D => n5765, CP => CLK_I, Q => 
                           n_2514, QN => n3118);
   KEY_EXPAN0_reg_22_18_inst : FD1 port map( D => n5764, CP => CLK_I, Q => 
                           n_2515, QN => n3117);
   KEY_EXPAN0_reg_21_18_inst : FD1 port map( D => n5763, CP => CLK_I, Q => 
                           n_2516, QN => n3120);
   KEY_EXPAN0_reg_20_18_inst : FD1 port map( D => n5762, CP => CLK_I, Q => 
                           n_2517, QN => n3119);
   KEY_EXPAN0_reg_19_18_inst : FD1 port map( D => n5761, CP => CLK_I, Q => 
                           n_2518, QN => n3122);
   KEY_EXPAN0_reg_18_18_inst : FD1 port map( D => n5760, CP => CLK_I, Q => 
                           n_2519, QN => n3121);
   KEY_EXPAN0_reg_17_18_inst : FD1 port map( D => n5759, CP => CLK_I, Q => 
                           n_2520, QN => n3124);
   KEY_EXPAN0_reg_16_18_inst : FD1 port map( D => n5758, CP => CLK_I, Q => 
                           n_2521, QN => n3123);
   KEY_EXPAN0_reg_15_18_inst : FD1 port map( D => n5757, CP => CLK_I, Q => 
                           n_2522, QN => n3110);
   KEY_EXPAN0_reg_14_18_inst : FD1 port map( D => n5756, CP => CLK_I, Q => 
                           n_2523, QN => n3109);
   KEY_EXPAN0_reg_13_18_inst : FD1 port map( D => n5755, CP => CLK_I, Q => 
                           n_2524, QN => n3112);
   KEY_EXPAN0_reg_12_18_inst : FD1 port map( D => n5754, CP => CLK_I, Q => 
                           n_2525, QN => n3111);
   KEY_EXPAN0_reg_11_18_inst : FD1 port map( D => n5753, CP => CLK_I, Q => 
                           n_2526, QN => n3114);
   KEY_EXPAN0_reg_10_18_inst : FD1 port map( D => n5752, CP => CLK_I, Q => 
                           n_2527, QN => n3113);
   KEY_EXPAN0_reg_9_18_inst : FD1 port map( D => n5751, CP => CLK_I, Q => 
                           n_2528, QN => n3116);
   KEY_EXPAN0_reg_8_18_inst : FD1 port map( D => n5750, CP => CLK_I, Q => 
                           n_2529, QN => n3115);
   KEY_EXPAN0_reg_7_18_inst : FD1 port map( D => n5749, CP => CLK_I, Q => 
                           n_2530, QN => n3102);
   KEY_EXPAN0_reg_6_18_inst : FD1 port map( D => n5748, CP => CLK_I, Q => 
                           n_2531, QN => n3101);
   KEY_EXPAN0_reg_5_18_inst : FD1 port map( D => n5747, CP => CLK_I, Q => 
                           n_2532, QN => n3104);
   KEY_EXPAN0_reg_4_18_inst : FD1 port map( D => n5746, CP => CLK_I, Q => 
                           n_2533, QN => n3103);
   KEY_EXPAN0_reg_3_18_inst : FD1 port map( D => n5745, CP => CLK_I, Q => 
                           n_2534, QN => n3106);
   KEY_EXPAN0_reg_2_18_inst : FD1 port map( D => n5744, CP => CLK_I, Q => 
                           n_2535, QN => n3105);
   KEY_EXPAN0_reg_1_18_inst : FD1 port map( D => n5743, CP => CLK_I, Q => 
                           n_2536, QN => n3108);
   KEY_EXPAN0_reg_0_18_inst : FD1 port map( D => n5742, CP => CLK_I, Q => 
                           n_2537, QN => n3107);
   v_KEY_COL_OUT0_reg_18_inst : FD1 port map( D => n4558, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_18_port, QN => n389);
   v_TEMP_VECTOR_reg_10_inst : FD1 port map( D => n6685, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_10_port, QN => n_2538);
   KEY_EXPAN0_reg_63_10_inst : FD1 port map( D => n5293, CP => CLK_I, Q => 
                           n_2539, QN => n3030);
   KEY_EXPAN0_reg_62_10_inst : FD1 port map( D => n5292, CP => CLK_I, Q => 
                           n_2540, QN => n3029);
   KEY_EXPAN0_reg_61_10_inst : FD1 port map( D => n5291, CP => CLK_I, Q => 
                           n_2541, QN => n3032);
   KEY_EXPAN0_reg_60_10_inst : FD1 port map( D => n5290, CP => CLK_I, Q => 
                           n_2542, QN => n3031);
   KEY_EXPAN0_reg_59_10_inst : FD1 port map( D => n5289, CP => CLK_I, Q => 
                           n_2543, QN => n3034);
   KEY_EXPAN0_reg_58_10_inst : FD1 port map( D => n5288, CP => CLK_I, Q => 
                           n_2544, QN => n3033);
   KEY_EXPAN0_reg_57_10_inst : FD1 port map( D => n5287, CP => CLK_I, Q => 
                           n_2545, QN => n3036);
   KEY_EXPAN0_reg_56_10_inst : FD1 port map( D => n5286, CP => CLK_I, Q => 
                           n_2546, QN => n3035);
   KEY_EXPAN0_reg_55_10_inst : FD1 port map( D => n5285, CP => CLK_I, Q => 
                           n_2547, QN => n3022);
   KEY_EXPAN0_reg_54_10_inst : FD1 port map( D => n5284, CP => CLK_I, Q => 
                           n_2548, QN => n3021);
   KEY_EXPAN0_reg_53_10_inst : FD1 port map( D => n5283, CP => CLK_I, Q => 
                           n_2549, QN => n3024);
   KEY_EXPAN0_reg_52_10_inst : FD1 port map( D => n5282, CP => CLK_I, Q => 
                           n_2550, QN => n3023);
   KEY_EXPAN0_reg_51_10_inst : FD1 port map( D => n5281, CP => CLK_I, Q => 
                           n_2551, QN => n3026);
   KEY_EXPAN0_reg_50_10_inst : FD1 port map( D => n5280, CP => CLK_I, Q => 
                           n_2552, QN => n3025);
   KEY_EXPAN0_reg_49_10_inst : FD1 port map( D => n5279, CP => CLK_I, Q => 
                           n_2553, QN => n3028);
   KEY_EXPAN0_reg_48_10_inst : FD1 port map( D => n5278, CP => CLK_I, Q => 
                           n_2554, QN => n3027);
   KEY_EXPAN0_reg_47_10_inst : FD1 port map( D => n5277, CP => CLK_I, Q => 
                           n_2555, QN => n3014);
   KEY_EXPAN0_reg_46_10_inst : FD1 port map( D => n5276, CP => CLK_I, Q => 
                           n_2556, QN => n3013);
   KEY_EXPAN0_reg_45_10_inst : FD1 port map( D => n5275, CP => CLK_I, Q => 
                           n_2557, QN => n3016);
   KEY_EXPAN0_reg_44_10_inst : FD1 port map( D => n5274, CP => CLK_I, Q => 
                           n_2558, QN => n3015);
   KEY_EXPAN0_reg_43_10_inst : FD1 port map( D => n5273, CP => CLK_I, Q => 
                           n_2559, QN => n3018);
   KEY_EXPAN0_reg_42_10_inst : FD1 port map( D => n5272, CP => CLK_I, Q => 
                           n_2560, QN => n3017);
   KEY_EXPAN0_reg_41_10_inst : FD1 port map( D => n5271, CP => CLK_I, Q => 
                           n_2561, QN => n3020);
   KEY_EXPAN0_reg_40_10_inst : FD1 port map( D => n5270, CP => CLK_I, Q => 
                           n_2562, QN => n3019);
   KEY_EXPAN0_reg_39_10_inst : FD1 port map( D => n5269, CP => CLK_I, Q => 
                           n_2563, QN => n3006);
   KEY_EXPAN0_reg_38_10_inst : FD1 port map( D => n5268, CP => CLK_I, Q => 
                           n_2564, QN => n3005);
   KEY_EXPAN0_reg_37_10_inst : FD1 port map( D => n5267, CP => CLK_I, Q => 
                           n_2565, QN => n3008);
   KEY_EXPAN0_reg_36_10_inst : FD1 port map( D => n5266, CP => CLK_I, Q => 
                           n_2566, QN => n3007);
   KEY_EXPAN0_reg_35_10_inst : FD1 port map( D => n5265, CP => CLK_I, Q => 
                           n_2567, QN => n3010);
   KEY_EXPAN0_reg_34_10_inst : FD1 port map( D => n5264, CP => CLK_I, Q => 
                           n_2568, QN => n3009);
   KEY_EXPAN0_reg_33_10_inst : FD1 port map( D => n5263, CP => CLK_I, Q => 
                           n_2569, QN => n3012);
   KEY_EXPAN0_reg_32_10_inst : FD1 port map( D => n5262, CP => CLK_I, Q => 
                           n_2570, QN => n3011);
   KEY_EXPAN0_reg_31_10_inst : FD1 port map( D => n5261, CP => CLK_I, Q => 
                           n_2571, QN => n3062);
   KEY_EXPAN0_reg_30_10_inst : FD1 port map( D => n5260, CP => CLK_I, Q => 
                           n_2572, QN => n3061);
   KEY_EXPAN0_reg_29_10_inst : FD1 port map( D => n5259, CP => CLK_I, Q => 
                           n_2573, QN => n3064);
   KEY_EXPAN0_reg_28_10_inst : FD1 port map( D => n5258, CP => CLK_I, Q => 
                           n_2574, QN => n3063);
   KEY_EXPAN0_reg_27_10_inst : FD1 port map( D => n5257, CP => CLK_I, Q => 
                           n_2575, QN => n3066);
   KEY_EXPAN0_reg_26_10_inst : FD1 port map( D => n5256, CP => CLK_I, Q => 
                           n_2576, QN => n3065);
   KEY_EXPAN0_reg_25_10_inst : FD1 port map( D => n5255, CP => CLK_I, Q => 
                           n_2577, QN => n3068);
   KEY_EXPAN0_reg_24_10_inst : FD1 port map( D => n5254, CP => CLK_I, Q => 
                           n_2578, QN => n3067);
   KEY_EXPAN0_reg_23_10_inst : FD1 port map( D => n5253, CP => CLK_I, Q => 
                           n_2579, QN => n3054);
   KEY_EXPAN0_reg_22_10_inst : FD1 port map( D => n5252, CP => CLK_I, Q => 
                           n_2580, QN => n3053);
   KEY_EXPAN0_reg_21_10_inst : FD1 port map( D => n5251, CP => CLK_I, Q => 
                           n_2581, QN => n3056);
   KEY_EXPAN0_reg_20_10_inst : FD1 port map( D => n5250, CP => CLK_I, Q => 
                           n_2582, QN => n3055);
   KEY_EXPAN0_reg_19_10_inst : FD1 port map( D => n5249, CP => CLK_I, Q => 
                           n_2583, QN => n3058);
   KEY_EXPAN0_reg_18_10_inst : FD1 port map( D => n5248, CP => CLK_I, Q => 
                           n_2584, QN => n3057);
   KEY_EXPAN0_reg_17_10_inst : FD1 port map( D => n5247, CP => CLK_I, Q => 
                           n_2585, QN => n3060);
   KEY_EXPAN0_reg_16_10_inst : FD1 port map( D => n5246, CP => CLK_I, Q => 
                           n_2586, QN => n3059);
   KEY_EXPAN0_reg_15_10_inst : FD1 port map( D => n5245, CP => CLK_I, Q => 
                           n_2587, QN => n3046);
   KEY_EXPAN0_reg_14_10_inst : FD1 port map( D => n5244, CP => CLK_I, Q => 
                           n_2588, QN => n3045);
   KEY_EXPAN0_reg_13_10_inst : FD1 port map( D => n5243, CP => CLK_I, Q => 
                           n_2589, QN => n3048);
   KEY_EXPAN0_reg_12_10_inst : FD1 port map( D => n5242, CP => CLK_I, Q => 
                           n_2590, QN => n3047);
   KEY_EXPAN0_reg_11_10_inst : FD1 port map( D => n5241, CP => CLK_I, Q => 
                           n_2591, QN => n3050);
   KEY_EXPAN0_reg_10_10_inst : FD1 port map( D => n5240, CP => CLK_I, Q => 
                           n_2592, QN => n3049);
   KEY_EXPAN0_reg_9_10_inst : FD1 port map( D => n5239, CP => CLK_I, Q => 
                           n_2593, QN => n3052);
   KEY_EXPAN0_reg_8_10_inst : FD1 port map( D => n5238, CP => CLK_I, Q => 
                           n_2594, QN => n3051);
   KEY_EXPAN0_reg_7_10_inst : FD1 port map( D => n5237, CP => CLK_I, Q => 
                           n_2595, QN => n3038);
   KEY_EXPAN0_reg_6_10_inst : FD1 port map( D => n5236, CP => CLK_I, Q => 
                           n_2596, QN => n3037);
   KEY_EXPAN0_reg_5_10_inst : FD1 port map( D => n5235, CP => CLK_I, Q => 
                           n_2597, QN => n3040);
   KEY_EXPAN0_reg_4_10_inst : FD1 port map( D => n5234, CP => CLK_I, Q => 
                           n_2598, QN => n3039);
   KEY_EXPAN0_reg_3_10_inst : FD1 port map( D => n5233, CP => CLK_I, Q => 
                           n_2599, QN => n3042);
   KEY_EXPAN0_reg_2_10_inst : FD1 port map( D => n5232, CP => CLK_I, Q => 
                           n_2600, QN => n3041);
   KEY_EXPAN0_reg_1_10_inst : FD1 port map( D => n5231, CP => CLK_I, Q => 
                           n_2601, QN => n3044);
   KEY_EXPAN0_reg_0_10_inst : FD1 port map( D => n5230, CP => CLK_I, Q => 
                           n_2602, QN => n3043);
   v_KEY_COL_OUT0_reg_10_inst : FD1 port map( D => n4557, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_10_port, QN => n327);
   v_TEMP_VECTOR_reg_1_inst : FD1 port map( D => n6694, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_1_port, QN => n_2603);
   KEY_EXPAN0_reg_63_1_inst : FD1 port map( D => n4717, CP => CLK_I, Q => 
                           n_2604, QN => n2966);
   KEY_EXPAN0_reg_62_1_inst : FD1 port map( D => n4716, CP => CLK_I, Q => 
                           n_2605, QN => n2965);
   KEY_EXPAN0_reg_61_1_inst : FD1 port map( D => n4715, CP => CLK_I, Q => 
                           n_2606, QN => n2968);
   KEY_EXPAN0_reg_60_1_inst : FD1 port map( D => n4714, CP => CLK_I, Q => 
                           n_2607, QN => n2967);
   KEY_EXPAN0_reg_59_1_inst : FD1 port map( D => n4713, CP => CLK_I, Q => 
                           n_2608, QN => n2970);
   KEY_EXPAN0_reg_58_1_inst : FD1 port map( D => n4712, CP => CLK_I, Q => 
                           n_2609, QN => n2969);
   KEY_EXPAN0_reg_57_1_inst : FD1 port map( D => n4711, CP => CLK_I, Q => 
                           n_2610, QN => n2972);
   KEY_EXPAN0_reg_56_1_inst : FD1 port map( D => n4710, CP => CLK_I, Q => 
                           n_2611, QN => n2971);
   KEY_EXPAN0_reg_55_1_inst : FD1 port map( D => n4709, CP => CLK_I, Q => 
                           n_2612, QN => n2958);
   KEY_EXPAN0_reg_54_1_inst : FD1 port map( D => n4708, CP => CLK_I, Q => 
                           n_2613, QN => n2957);
   KEY_EXPAN0_reg_53_1_inst : FD1 port map( D => n4707, CP => CLK_I, Q => 
                           n_2614, QN => n2960);
   KEY_EXPAN0_reg_52_1_inst : FD1 port map( D => n4706, CP => CLK_I, Q => 
                           n_2615, QN => n2959);
   KEY_EXPAN0_reg_51_1_inst : FD1 port map( D => n4705, CP => CLK_I, Q => 
                           n_2616, QN => n2962);
   KEY_EXPAN0_reg_50_1_inst : FD1 port map( D => n4704, CP => CLK_I, Q => 
                           n_2617, QN => n2961);
   KEY_EXPAN0_reg_49_1_inst : FD1 port map( D => n4703, CP => CLK_I, Q => 
                           n_2618, QN => n2964);
   KEY_EXPAN0_reg_48_1_inst : FD1 port map( D => n4702, CP => CLK_I, Q => 
                           n_2619, QN => n2963);
   KEY_EXPAN0_reg_47_1_inst : FD1 port map( D => n4701, CP => CLK_I, Q => 
                           n_2620, QN => n2950);
   KEY_EXPAN0_reg_46_1_inst : FD1 port map( D => n4700, CP => CLK_I, Q => 
                           n_2621, QN => n2949);
   KEY_EXPAN0_reg_45_1_inst : FD1 port map( D => n4699, CP => CLK_I, Q => 
                           n_2622, QN => n2952);
   KEY_EXPAN0_reg_44_1_inst : FD1 port map( D => n4698, CP => CLK_I, Q => 
                           n_2623, QN => n2951);
   KEY_EXPAN0_reg_43_1_inst : FD1 port map( D => n4697, CP => CLK_I, Q => 
                           n_2624, QN => n2954);
   KEY_EXPAN0_reg_42_1_inst : FD1 port map( D => n4696, CP => CLK_I, Q => 
                           n_2625, QN => n2953);
   KEY_EXPAN0_reg_41_1_inst : FD1 port map( D => n4695, CP => CLK_I, Q => 
                           n_2626, QN => n2956);
   KEY_EXPAN0_reg_40_1_inst : FD1 port map( D => n4694, CP => CLK_I, Q => 
                           n_2627, QN => n2955);
   KEY_EXPAN0_reg_39_1_inst : FD1 port map( D => n4693, CP => CLK_I, Q => 
                           n_2628, QN => n2942);
   KEY_EXPAN0_reg_38_1_inst : FD1 port map( D => n4692, CP => CLK_I, Q => 
                           n_2629, QN => n2941);
   KEY_EXPAN0_reg_37_1_inst : FD1 port map( D => n4691, CP => CLK_I, Q => 
                           n_2630, QN => n2944);
   KEY_EXPAN0_reg_36_1_inst : FD1 port map( D => n4690, CP => CLK_I, Q => 
                           n_2631, QN => n2943);
   KEY_EXPAN0_reg_35_1_inst : FD1 port map( D => n4689, CP => CLK_I, Q => 
                           n_2632, QN => n2946);
   KEY_EXPAN0_reg_34_1_inst : FD1 port map( D => n4688, CP => CLK_I, Q => 
                           n_2633, QN => n2945);
   KEY_EXPAN0_reg_33_1_inst : FD1 port map( D => n4687, CP => CLK_I, Q => 
                           n_2634, QN => n2948);
   KEY_EXPAN0_reg_32_1_inst : FD1 port map( D => n4686, CP => CLK_I, Q => 
                           n_2635, QN => n2947);
   KEY_EXPAN0_reg_31_1_inst : FD1 port map( D => n4685, CP => CLK_I, Q => 
                           n_2636, QN => n2998);
   KEY_EXPAN0_reg_30_1_inst : FD1 port map( D => n4684, CP => CLK_I, Q => 
                           n_2637, QN => n2997);
   KEY_EXPAN0_reg_29_1_inst : FD1 port map( D => n4683, CP => CLK_I, Q => 
                           n_2638, QN => n3000);
   KEY_EXPAN0_reg_28_1_inst : FD1 port map( D => n4682, CP => CLK_I, Q => 
                           n_2639, QN => n2999);
   KEY_EXPAN0_reg_27_1_inst : FD1 port map( D => n4681, CP => CLK_I, Q => 
                           n_2640, QN => n3002);
   KEY_EXPAN0_reg_26_1_inst : FD1 port map( D => n4680, CP => CLK_I, Q => 
                           n_2641, QN => n3001);
   KEY_EXPAN0_reg_25_1_inst : FD1 port map( D => n4679, CP => CLK_I, Q => 
                           n_2642, QN => n3004);
   KEY_EXPAN0_reg_24_1_inst : FD1 port map( D => n4678, CP => CLK_I, Q => 
                           n_2643, QN => n3003);
   KEY_EXPAN0_reg_23_1_inst : FD1 port map( D => n4677, CP => CLK_I, Q => 
                           n_2644, QN => n2990);
   KEY_EXPAN0_reg_22_1_inst : FD1 port map( D => n4676, CP => CLK_I, Q => 
                           n_2645, QN => n2989);
   KEY_EXPAN0_reg_21_1_inst : FD1 port map( D => n4675, CP => CLK_I, Q => 
                           n_2646, QN => n2992);
   KEY_EXPAN0_reg_20_1_inst : FD1 port map( D => n4674, CP => CLK_I, Q => 
                           n_2647, QN => n2991);
   KEY_EXPAN0_reg_19_1_inst : FD1 port map( D => n4673, CP => CLK_I, Q => 
                           n_2648, QN => n2994);
   KEY_EXPAN0_reg_18_1_inst : FD1 port map( D => n4672, CP => CLK_I, Q => 
                           n_2649, QN => n2993);
   KEY_EXPAN0_reg_17_1_inst : FD1 port map( D => n4671, CP => CLK_I, Q => 
                           n_2650, QN => n2996);
   KEY_EXPAN0_reg_16_1_inst : FD1 port map( D => n4670, CP => CLK_I, Q => 
                           n_2651, QN => n2995);
   KEY_EXPAN0_reg_15_1_inst : FD1 port map( D => n4669, CP => CLK_I, Q => 
                           n_2652, QN => n2982);
   KEY_EXPAN0_reg_14_1_inst : FD1 port map( D => n4668, CP => CLK_I, Q => 
                           n_2653, QN => n2981);
   KEY_EXPAN0_reg_13_1_inst : FD1 port map( D => n4667, CP => CLK_I, Q => 
                           n_2654, QN => n2984);
   KEY_EXPAN0_reg_12_1_inst : FD1 port map( D => n4666, CP => CLK_I, Q => 
                           n_2655, QN => n2983);
   KEY_EXPAN0_reg_11_1_inst : FD1 port map( D => n4665, CP => CLK_I, Q => 
                           n_2656, QN => n2986);
   KEY_EXPAN0_reg_10_1_inst : FD1 port map( D => n4664, CP => CLK_I, Q => 
                           n_2657, QN => n2985);
   KEY_EXPAN0_reg_9_1_inst : FD1 port map( D => n4663, CP => CLK_I, Q => n_2658
                           , QN => n2988);
   KEY_EXPAN0_reg_8_1_inst : FD1 port map( D => n4662, CP => CLK_I, Q => n_2659
                           , QN => n2987);
   KEY_EXPAN0_reg_7_1_inst : FD1 port map( D => n4661, CP => CLK_I, Q => n_2660
                           , QN => n2974);
   KEY_EXPAN0_reg_6_1_inst : FD1 port map( D => n4660, CP => CLK_I, Q => n_2661
                           , QN => n2973);
   KEY_EXPAN0_reg_5_1_inst : FD1 port map( D => n4659, CP => CLK_I, Q => n_2662
                           , QN => n2976);
   KEY_EXPAN0_reg_4_1_inst : FD1 port map( D => n4658, CP => CLK_I, Q => n_2663
                           , QN => n2975);
   KEY_EXPAN0_reg_3_1_inst : FD1 port map( D => n4657, CP => CLK_I, Q => n_2664
                           , QN => n2978);
   KEY_EXPAN0_reg_2_1_inst : FD1 port map( D => n4656, CP => CLK_I, Q => n_2665
                           , QN => n2977);
   KEY_EXPAN0_reg_1_1_inst : FD1 port map( D => n4655, CP => CLK_I, Q => n_2666
                           , QN => n2980);
   KEY_EXPAN0_reg_0_1_inst : FD1 port map( D => n4654, CP => CLK_I, Q => n_2667
                           , QN => n2979);
   v_KEY_COL_OUT0_reg_1_inst : FD1 port map( D => n4556, CP => CLK_I, Q => 
                           n_2668, QN => n1542);
   v_TEMP_VECTOR_reg_25_inst : FD1 port map( D => n6670, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_25_port, QN => n_2669);
   KEY_EXPAN0_reg_63_25_inst : FD1 port map( D => n6253, CP => CLK_I, Q => 
                           n_2670, QN => n2902);
   KEY_EXPAN0_reg_62_25_inst : FD1 port map( D => n6252, CP => CLK_I, Q => 
                           n_2671, QN => n2901);
   KEY_EXPAN0_reg_61_25_inst : FD1 port map( D => n6251, CP => CLK_I, Q => 
                           n_2672, QN => n2904);
   KEY_EXPAN0_reg_60_25_inst : FD1 port map( D => n6250, CP => CLK_I, Q => 
                           n_2673, QN => n2903);
   KEY_EXPAN0_reg_59_25_inst : FD1 port map( D => n6249, CP => CLK_I, Q => 
                           n_2674, QN => n2906);
   KEY_EXPAN0_reg_58_25_inst : FD1 port map( D => n6248, CP => CLK_I, Q => 
                           n_2675, QN => n2905);
   KEY_EXPAN0_reg_57_25_inst : FD1 port map( D => n6247, CP => CLK_I, Q => 
                           n_2676, QN => n2908);
   KEY_EXPAN0_reg_56_25_inst : FD1 port map( D => n6246, CP => CLK_I, Q => 
                           n_2677, QN => n2907);
   KEY_EXPAN0_reg_55_25_inst : FD1 port map( D => n6245, CP => CLK_I, Q => 
                           n_2678, QN => n2894);
   KEY_EXPAN0_reg_54_25_inst : FD1 port map( D => n6244, CP => CLK_I, Q => 
                           n_2679, QN => n2893);
   KEY_EXPAN0_reg_53_25_inst : FD1 port map( D => n6243, CP => CLK_I, Q => 
                           n_2680, QN => n2896);
   KEY_EXPAN0_reg_52_25_inst : FD1 port map( D => n6242, CP => CLK_I, Q => 
                           n_2681, QN => n2895);
   KEY_EXPAN0_reg_51_25_inst : FD1 port map( D => n6241, CP => CLK_I, Q => 
                           n_2682, QN => n2898);
   KEY_EXPAN0_reg_50_25_inst : FD1 port map( D => n6240, CP => CLK_I, Q => 
                           n_2683, QN => n2897);
   KEY_EXPAN0_reg_49_25_inst : FD1 port map( D => n6239, CP => CLK_I, Q => 
                           n_2684, QN => n2900);
   KEY_EXPAN0_reg_48_25_inst : FD1 port map( D => n6238, CP => CLK_I, Q => 
                           n_2685, QN => n2899);
   KEY_EXPAN0_reg_47_25_inst : FD1 port map( D => n6237, CP => CLK_I, Q => 
                           n_2686, QN => n2886);
   KEY_EXPAN0_reg_46_25_inst : FD1 port map( D => n6236, CP => CLK_I, Q => 
                           n_2687, QN => n2885);
   KEY_EXPAN0_reg_45_25_inst : FD1 port map( D => n6235, CP => CLK_I, Q => 
                           n_2688, QN => n2888);
   KEY_EXPAN0_reg_44_25_inst : FD1 port map( D => n6234, CP => CLK_I, Q => 
                           n_2689, QN => n2887);
   KEY_EXPAN0_reg_43_25_inst : FD1 port map( D => n6233, CP => CLK_I, Q => 
                           n_2690, QN => n2890);
   KEY_EXPAN0_reg_42_25_inst : FD1 port map( D => n6232, CP => CLK_I, Q => 
                           n_2691, QN => n2889);
   KEY_EXPAN0_reg_41_25_inst : FD1 port map( D => n6231, CP => CLK_I, Q => 
                           n_2692, QN => n2892);
   KEY_EXPAN0_reg_40_25_inst : FD1 port map( D => n6230, CP => CLK_I, Q => 
                           n_2693, QN => n2891);
   KEY_EXPAN0_reg_39_25_inst : FD1 port map( D => n6229, CP => CLK_I, Q => 
                           n_2694, QN => n2878);
   KEY_EXPAN0_reg_38_25_inst : FD1 port map( D => n6228, CP => CLK_I, Q => 
                           n_2695, QN => n2877);
   KEY_EXPAN0_reg_37_25_inst : FD1 port map( D => n6227, CP => CLK_I, Q => 
                           n_2696, QN => n2880);
   KEY_EXPAN0_reg_36_25_inst : FD1 port map( D => n6226, CP => CLK_I, Q => 
                           n_2697, QN => n2879);
   KEY_EXPAN0_reg_35_25_inst : FD1 port map( D => n6225, CP => CLK_I, Q => 
                           n_2698, QN => n2882);
   KEY_EXPAN0_reg_34_25_inst : FD1 port map( D => n6224, CP => CLK_I, Q => 
                           n_2699, QN => n2881);
   KEY_EXPAN0_reg_33_25_inst : FD1 port map( D => n6223, CP => CLK_I, Q => 
                           n_2700, QN => n2884);
   KEY_EXPAN0_reg_32_25_inst : FD1 port map( D => n6222, CP => CLK_I, Q => 
                           n_2701, QN => n2883);
   KEY_EXPAN0_reg_31_25_inst : FD1 port map( D => n6221, CP => CLK_I, Q => 
                           n_2702, QN => n2934);
   KEY_EXPAN0_reg_30_25_inst : FD1 port map( D => n6220, CP => CLK_I, Q => 
                           n_2703, QN => n2933);
   KEY_EXPAN0_reg_29_25_inst : FD1 port map( D => n6219, CP => CLK_I, Q => 
                           n_2704, QN => n2936);
   KEY_EXPAN0_reg_28_25_inst : FD1 port map( D => n6218, CP => CLK_I, Q => 
                           n_2705, QN => n2935);
   KEY_EXPAN0_reg_27_25_inst : FD1 port map( D => n6217, CP => CLK_I, Q => 
                           n_2706, QN => n2938);
   KEY_EXPAN0_reg_26_25_inst : FD1 port map( D => n6216, CP => CLK_I, Q => 
                           n_2707, QN => n2937);
   KEY_EXPAN0_reg_25_25_inst : FD1 port map( D => n6215, CP => CLK_I, Q => 
                           n_2708, QN => n2940);
   KEY_EXPAN0_reg_24_25_inst : FD1 port map( D => n6214, CP => CLK_I, Q => 
                           n_2709, QN => n2939);
   KEY_EXPAN0_reg_23_25_inst : FD1 port map( D => n6213, CP => CLK_I, Q => 
                           n_2710, QN => n2926);
   KEY_EXPAN0_reg_22_25_inst : FD1 port map( D => n6212, CP => CLK_I, Q => 
                           n_2711, QN => n2925);
   KEY_EXPAN0_reg_21_25_inst : FD1 port map( D => n6211, CP => CLK_I, Q => 
                           n_2712, QN => n2928);
   KEY_EXPAN0_reg_20_25_inst : FD1 port map( D => n6210, CP => CLK_I, Q => 
                           n_2713, QN => n2927);
   KEY_EXPAN0_reg_19_25_inst : FD1 port map( D => n6209, CP => CLK_I, Q => 
                           n_2714, QN => n2930);
   KEY_EXPAN0_reg_18_25_inst : FD1 port map( D => n6208, CP => CLK_I, Q => 
                           n_2715, QN => n2929);
   KEY_EXPAN0_reg_17_25_inst : FD1 port map( D => n6207, CP => CLK_I, Q => 
                           n_2716, QN => n2932);
   KEY_EXPAN0_reg_16_25_inst : FD1 port map( D => n6206, CP => CLK_I, Q => 
                           n_2717, QN => n2931);
   KEY_EXPAN0_reg_15_25_inst : FD1 port map( D => n6205, CP => CLK_I, Q => 
                           n_2718, QN => n2918);
   KEY_EXPAN0_reg_14_25_inst : FD1 port map( D => n6204, CP => CLK_I, Q => 
                           n_2719, QN => n2917);
   KEY_EXPAN0_reg_13_25_inst : FD1 port map( D => n6203, CP => CLK_I, Q => 
                           n_2720, QN => n2920);
   KEY_EXPAN0_reg_12_25_inst : FD1 port map( D => n6202, CP => CLK_I, Q => 
                           n_2721, QN => n2919);
   KEY_EXPAN0_reg_11_25_inst : FD1 port map( D => n6201, CP => CLK_I, Q => 
                           n_2722, QN => n2922);
   KEY_EXPAN0_reg_10_25_inst : FD1 port map( D => n6200, CP => CLK_I, Q => 
                           n_2723, QN => n2921);
   KEY_EXPAN0_reg_9_25_inst : FD1 port map( D => n6199, CP => CLK_I, Q => 
                           n_2724, QN => n2924);
   KEY_EXPAN0_reg_8_25_inst : FD1 port map( D => n6198, CP => CLK_I, Q => 
                           n_2725, QN => n2923);
   KEY_EXPAN0_reg_7_25_inst : FD1 port map( D => n6197, CP => CLK_I, Q => 
                           n_2726, QN => n2910);
   KEY_EXPAN0_reg_6_25_inst : FD1 port map( D => n6196, CP => CLK_I, Q => 
                           n_2727, QN => n2909);
   KEY_EXPAN0_reg_5_25_inst : FD1 port map( D => n6195, CP => CLK_I, Q => 
                           n_2728, QN => n2912);
   KEY_EXPAN0_reg_4_25_inst : FD1 port map( D => n6194, CP => CLK_I, Q => 
                           n_2729, QN => n2911);
   KEY_EXPAN0_reg_3_25_inst : FD1 port map( D => n6193, CP => CLK_I, Q => 
                           n_2730, QN => n2914);
   KEY_EXPAN0_reg_2_25_inst : FD1 port map( D => n6192, CP => CLK_I, Q => 
                           n_2731, QN => n2913);
   KEY_EXPAN0_reg_1_25_inst : FD1 port map( D => n6191, CP => CLK_I, Q => 
                           n_2732, QN => n2916);
   KEY_EXPAN0_reg_0_25_inst : FD1 port map( D => n6190, CP => CLK_I, Q => 
                           n_2733, QN => n2915);
   v_KEY_COL_OUT0_reg_25_inst : FD1 port map( D => n4555, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_25_port, QN => n1454);
   v_TEMP_VECTOR_reg_17_inst : FD1 port map( D => n6678, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_17_port, QN => n_2734);
   KEY_EXPAN0_reg_63_17_inst : FD1 port map( D => n5741, CP => CLK_I, Q => 
                           n_2735, QN => n2838);
   KEY_EXPAN0_reg_62_17_inst : FD1 port map( D => n5740, CP => CLK_I, Q => 
                           n_2736, QN => n2837);
   KEY_EXPAN0_reg_61_17_inst : FD1 port map( D => n5739, CP => CLK_I, Q => 
                           n_2737, QN => n2840);
   KEY_EXPAN0_reg_60_17_inst : FD1 port map( D => n5738, CP => CLK_I, Q => 
                           n_2738, QN => n2839);
   KEY_EXPAN0_reg_59_17_inst : FD1 port map( D => n5737, CP => CLK_I, Q => 
                           n_2739, QN => n2842);
   KEY_EXPAN0_reg_58_17_inst : FD1 port map( D => n5736, CP => CLK_I, Q => 
                           n_2740, QN => n2841);
   KEY_EXPAN0_reg_57_17_inst : FD1 port map( D => n5735, CP => CLK_I, Q => 
                           n_2741, QN => n2844);
   KEY_EXPAN0_reg_56_17_inst : FD1 port map( D => n5734, CP => CLK_I, Q => 
                           n_2742, QN => n2843);
   KEY_EXPAN0_reg_55_17_inst : FD1 port map( D => n5733, CP => CLK_I, Q => 
                           n_2743, QN => n2830);
   KEY_EXPAN0_reg_54_17_inst : FD1 port map( D => n5732, CP => CLK_I, Q => 
                           n_2744, QN => n2829);
   KEY_EXPAN0_reg_53_17_inst : FD1 port map( D => n5731, CP => CLK_I, Q => 
                           n_2745, QN => n2832);
   KEY_EXPAN0_reg_52_17_inst : FD1 port map( D => n5730, CP => CLK_I, Q => 
                           n_2746, QN => n2831);
   KEY_EXPAN0_reg_51_17_inst : FD1 port map( D => n5729, CP => CLK_I, Q => 
                           n_2747, QN => n2834);
   KEY_EXPAN0_reg_50_17_inst : FD1 port map( D => n5728, CP => CLK_I, Q => 
                           n_2748, QN => n2833);
   KEY_EXPAN0_reg_49_17_inst : FD1 port map( D => n5727, CP => CLK_I, Q => 
                           n_2749, QN => n2836);
   KEY_EXPAN0_reg_48_17_inst : FD1 port map( D => n5726, CP => CLK_I, Q => 
                           n_2750, QN => n2835);
   KEY_EXPAN0_reg_47_17_inst : FD1 port map( D => n5725, CP => CLK_I, Q => 
                           n_2751, QN => n2822);
   KEY_EXPAN0_reg_46_17_inst : FD1 port map( D => n5724, CP => CLK_I, Q => 
                           n_2752, QN => n2821);
   KEY_EXPAN0_reg_45_17_inst : FD1 port map( D => n5723, CP => CLK_I, Q => 
                           n_2753, QN => n2824);
   KEY_EXPAN0_reg_44_17_inst : FD1 port map( D => n5722, CP => CLK_I, Q => 
                           n_2754, QN => n2823);
   KEY_EXPAN0_reg_43_17_inst : FD1 port map( D => n5721, CP => CLK_I, Q => 
                           n_2755, QN => n2826);
   KEY_EXPAN0_reg_42_17_inst : FD1 port map( D => n5720, CP => CLK_I, Q => 
                           n_2756, QN => n2825);
   KEY_EXPAN0_reg_41_17_inst : FD1 port map( D => n5719, CP => CLK_I, Q => 
                           n_2757, QN => n2828);
   KEY_EXPAN0_reg_40_17_inst : FD1 port map( D => n5718, CP => CLK_I, Q => 
                           n_2758, QN => n2827);
   KEY_EXPAN0_reg_39_17_inst : FD1 port map( D => n5717, CP => CLK_I, Q => 
                           n_2759, QN => n2814);
   KEY_EXPAN0_reg_38_17_inst : FD1 port map( D => n5716, CP => CLK_I, Q => 
                           n_2760, QN => n2813);
   KEY_EXPAN0_reg_37_17_inst : FD1 port map( D => n5715, CP => CLK_I, Q => 
                           n_2761, QN => n2816);
   KEY_EXPAN0_reg_36_17_inst : FD1 port map( D => n5714, CP => CLK_I, Q => 
                           n_2762, QN => n2815);
   KEY_EXPAN0_reg_35_17_inst : FD1 port map( D => n5713, CP => CLK_I, Q => 
                           n_2763, QN => n2818);
   KEY_EXPAN0_reg_34_17_inst : FD1 port map( D => n5712, CP => CLK_I, Q => 
                           n_2764, QN => n2817);
   KEY_EXPAN0_reg_33_17_inst : FD1 port map( D => n5711, CP => CLK_I, Q => 
                           n_2765, QN => n2820);
   KEY_EXPAN0_reg_32_17_inst : FD1 port map( D => n5710, CP => CLK_I, Q => 
                           n_2766, QN => n2819);
   KEY_EXPAN0_reg_31_17_inst : FD1 port map( D => n5709, CP => CLK_I, Q => 
                           n_2767, QN => n2870);
   KEY_EXPAN0_reg_30_17_inst : FD1 port map( D => n5708, CP => CLK_I, Q => 
                           n_2768, QN => n2869);
   KEY_EXPAN0_reg_29_17_inst : FD1 port map( D => n5707, CP => CLK_I, Q => 
                           n_2769, QN => n2872);
   KEY_EXPAN0_reg_28_17_inst : FD1 port map( D => n5706, CP => CLK_I, Q => 
                           n_2770, QN => n2871);
   KEY_EXPAN0_reg_27_17_inst : FD1 port map( D => n5705, CP => CLK_I, Q => 
                           n_2771, QN => n2874);
   KEY_EXPAN0_reg_26_17_inst : FD1 port map( D => n5704, CP => CLK_I, Q => 
                           n_2772, QN => n2873);
   KEY_EXPAN0_reg_25_17_inst : FD1 port map( D => n5703, CP => CLK_I, Q => 
                           n_2773, QN => n2876);
   KEY_EXPAN0_reg_24_17_inst : FD1 port map( D => n5702, CP => CLK_I, Q => 
                           n_2774, QN => n2875);
   KEY_EXPAN0_reg_23_17_inst : FD1 port map( D => n5701, CP => CLK_I, Q => 
                           n_2775, QN => n2862);
   KEY_EXPAN0_reg_22_17_inst : FD1 port map( D => n5700, CP => CLK_I, Q => 
                           n_2776, QN => n2861);
   KEY_EXPAN0_reg_21_17_inst : FD1 port map( D => n5699, CP => CLK_I, Q => 
                           n_2777, QN => n2864);
   KEY_EXPAN0_reg_20_17_inst : FD1 port map( D => n5698, CP => CLK_I, Q => 
                           n_2778, QN => n2863);
   KEY_EXPAN0_reg_19_17_inst : FD1 port map( D => n5697, CP => CLK_I, Q => 
                           n_2779, QN => n2866);
   KEY_EXPAN0_reg_18_17_inst : FD1 port map( D => n5696, CP => CLK_I, Q => 
                           n_2780, QN => n2865);
   KEY_EXPAN0_reg_17_17_inst : FD1 port map( D => n5695, CP => CLK_I, Q => 
                           n_2781, QN => n2868);
   KEY_EXPAN0_reg_16_17_inst : FD1 port map( D => n5694, CP => CLK_I, Q => 
                           n_2782, QN => n2867);
   KEY_EXPAN0_reg_15_17_inst : FD1 port map( D => n5693, CP => CLK_I, Q => 
                           n_2783, QN => n2854);
   KEY_EXPAN0_reg_14_17_inst : FD1 port map( D => n5692, CP => CLK_I, Q => 
                           n_2784, QN => n2853);
   KEY_EXPAN0_reg_13_17_inst : FD1 port map( D => n5691, CP => CLK_I, Q => 
                           n_2785, QN => n2856);
   KEY_EXPAN0_reg_12_17_inst : FD1 port map( D => n5690, CP => CLK_I, Q => 
                           n_2786, QN => n2855);
   KEY_EXPAN0_reg_11_17_inst : FD1 port map( D => n5689, CP => CLK_I, Q => 
                           n_2787, QN => n2858);
   KEY_EXPAN0_reg_10_17_inst : FD1 port map( D => n5688, CP => CLK_I, Q => 
                           n_2788, QN => n2857);
   KEY_EXPAN0_reg_9_17_inst : FD1 port map( D => n5687, CP => CLK_I, Q => 
                           n_2789, QN => n2860);
   KEY_EXPAN0_reg_8_17_inst : FD1 port map( D => n5686, CP => CLK_I, Q => 
                           n_2790, QN => n2859);
   KEY_EXPAN0_reg_7_17_inst : FD1 port map( D => n5685, CP => CLK_I, Q => 
                           n_2791, QN => n2846);
   KEY_EXPAN0_reg_6_17_inst : FD1 port map( D => n5684, CP => CLK_I, Q => 
                           n_2792, QN => n2845);
   KEY_EXPAN0_reg_5_17_inst : FD1 port map( D => n5683, CP => CLK_I, Q => 
                           n_2793, QN => n2848);
   KEY_EXPAN0_reg_4_17_inst : FD1 port map( D => n5682, CP => CLK_I, Q => 
                           n_2794, QN => n2847);
   KEY_EXPAN0_reg_3_17_inst : FD1 port map( D => n5681, CP => CLK_I, Q => 
                           n_2795, QN => n2850);
   KEY_EXPAN0_reg_2_17_inst : FD1 port map( D => n5680, CP => CLK_I, Q => 
                           n_2796, QN => n2849);
   KEY_EXPAN0_reg_1_17_inst : FD1 port map( D => n5679, CP => CLK_I, Q => 
                           n_2797, QN => n2852);
   KEY_EXPAN0_reg_0_17_inst : FD1 port map( D => n5678, CP => CLK_I, Q => 
                           n_2798, QN => n2851);
   v_KEY_COL_OUT0_reg_17_inst : FD1 port map( D => n4554, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_17_port, QN => n1889);
   v_TEMP_VECTOR_reg_9_inst : FD1 port map( D => n6686, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_9_port, QN => n_2799);
   KEY_EXPAN0_reg_63_9_inst : FD1 port map( D => n5229, CP => CLK_I, Q => 
                           n_2800, QN => n2774);
   KEY_EXPAN0_reg_62_9_inst : FD1 port map( D => n5228, CP => CLK_I, Q => 
                           n_2801, QN => n2773);
   KEY_EXPAN0_reg_61_9_inst : FD1 port map( D => n5227, CP => CLK_I, Q => 
                           n_2802, QN => n2776);
   KEY_EXPAN0_reg_60_9_inst : FD1 port map( D => n5226, CP => CLK_I, Q => 
                           n_2803, QN => n2775);
   KEY_EXPAN0_reg_59_9_inst : FD1 port map( D => n5225, CP => CLK_I, Q => 
                           n_2804, QN => n2778);
   KEY_EXPAN0_reg_58_9_inst : FD1 port map( D => n5224, CP => CLK_I, Q => 
                           n_2805, QN => n2777);
   KEY_EXPAN0_reg_57_9_inst : FD1 port map( D => n5223, CP => CLK_I, Q => 
                           n_2806, QN => n2780);
   KEY_EXPAN0_reg_56_9_inst : FD1 port map( D => n5222, CP => CLK_I, Q => 
                           n_2807, QN => n2779);
   KEY_EXPAN0_reg_55_9_inst : FD1 port map( D => n5221, CP => CLK_I, Q => 
                           n_2808, QN => n2766);
   KEY_EXPAN0_reg_54_9_inst : FD1 port map( D => n5220, CP => CLK_I, Q => 
                           n_2809, QN => n2765);
   KEY_EXPAN0_reg_53_9_inst : FD1 port map( D => n5219, CP => CLK_I, Q => 
                           n_2810, QN => n2768);
   KEY_EXPAN0_reg_52_9_inst : FD1 port map( D => n5218, CP => CLK_I, Q => 
                           n_2811, QN => n2767);
   KEY_EXPAN0_reg_51_9_inst : FD1 port map( D => n5217, CP => CLK_I, Q => 
                           n_2812, QN => n2770);
   KEY_EXPAN0_reg_50_9_inst : FD1 port map( D => n5216, CP => CLK_I, Q => 
                           n_2813, QN => n2769);
   KEY_EXPAN0_reg_49_9_inst : FD1 port map( D => n5215, CP => CLK_I, Q => 
                           n_2814, QN => n2772);
   KEY_EXPAN0_reg_48_9_inst : FD1 port map( D => n5214, CP => CLK_I, Q => 
                           n_2815, QN => n2771);
   KEY_EXPAN0_reg_47_9_inst : FD1 port map( D => n5213, CP => CLK_I, Q => 
                           n_2816, QN => n2758);
   KEY_EXPAN0_reg_46_9_inst : FD1 port map( D => n5212, CP => CLK_I, Q => 
                           n_2817, QN => n2757);
   KEY_EXPAN0_reg_45_9_inst : FD1 port map( D => n5211, CP => CLK_I, Q => 
                           n_2818, QN => n2760);
   KEY_EXPAN0_reg_44_9_inst : FD1 port map( D => n5210, CP => CLK_I, Q => 
                           n_2819, QN => n2759);
   KEY_EXPAN0_reg_43_9_inst : FD1 port map( D => n5209, CP => CLK_I, Q => 
                           n_2820, QN => n2762);
   KEY_EXPAN0_reg_42_9_inst : FD1 port map( D => n5208, CP => CLK_I, Q => 
                           n_2821, QN => n2761);
   KEY_EXPAN0_reg_41_9_inst : FD1 port map( D => n5207, CP => CLK_I, Q => 
                           n_2822, QN => n2764);
   KEY_EXPAN0_reg_40_9_inst : FD1 port map( D => n5206, CP => CLK_I, Q => 
                           n_2823, QN => n2763);
   KEY_EXPAN0_reg_39_9_inst : FD1 port map( D => n5205, CP => CLK_I, Q => 
                           n_2824, QN => n2750);
   KEY_EXPAN0_reg_38_9_inst : FD1 port map( D => n5204, CP => CLK_I, Q => 
                           n_2825, QN => n2749);
   KEY_EXPAN0_reg_37_9_inst : FD1 port map( D => n5203, CP => CLK_I, Q => 
                           n_2826, QN => n2752);
   KEY_EXPAN0_reg_36_9_inst : FD1 port map( D => n5202, CP => CLK_I, Q => 
                           n_2827, QN => n2751);
   KEY_EXPAN0_reg_35_9_inst : FD1 port map( D => n5201, CP => CLK_I, Q => 
                           n_2828, QN => n2754);
   KEY_EXPAN0_reg_34_9_inst : FD1 port map( D => n5200, CP => CLK_I, Q => 
                           n_2829, QN => n2753);
   KEY_EXPAN0_reg_33_9_inst : FD1 port map( D => n5199, CP => CLK_I, Q => 
                           n_2830, QN => n2756);
   KEY_EXPAN0_reg_32_9_inst : FD1 port map( D => n5198, CP => CLK_I, Q => 
                           n_2831, QN => n2755);
   KEY_EXPAN0_reg_31_9_inst : FD1 port map( D => n5197, CP => CLK_I, Q => 
                           n_2832, QN => n2806);
   KEY_EXPAN0_reg_30_9_inst : FD1 port map( D => n5196, CP => CLK_I, Q => 
                           n_2833, QN => n2805);
   KEY_EXPAN0_reg_29_9_inst : FD1 port map( D => n5195, CP => CLK_I, Q => 
                           n_2834, QN => n2808);
   KEY_EXPAN0_reg_28_9_inst : FD1 port map( D => n5194, CP => CLK_I, Q => 
                           n_2835, QN => n2807);
   KEY_EXPAN0_reg_27_9_inst : FD1 port map( D => n5193, CP => CLK_I, Q => 
                           n_2836, QN => n2810);
   KEY_EXPAN0_reg_26_9_inst : FD1 port map( D => n5192, CP => CLK_I, Q => 
                           n_2837, QN => n2809);
   KEY_EXPAN0_reg_25_9_inst : FD1 port map( D => n5191, CP => CLK_I, Q => 
                           n_2838, QN => n2812);
   KEY_EXPAN0_reg_24_9_inst : FD1 port map( D => n5190, CP => CLK_I, Q => 
                           n_2839, QN => n2811);
   KEY_EXPAN0_reg_23_9_inst : FD1 port map( D => n5189, CP => CLK_I, Q => 
                           n_2840, QN => n2798);
   KEY_EXPAN0_reg_22_9_inst : FD1 port map( D => n5188, CP => CLK_I, Q => 
                           n_2841, QN => n2797);
   KEY_EXPAN0_reg_21_9_inst : FD1 port map( D => n5187, CP => CLK_I, Q => 
                           n_2842, QN => n2800);
   KEY_EXPAN0_reg_20_9_inst : FD1 port map( D => n5186, CP => CLK_I, Q => 
                           n_2843, QN => n2799);
   KEY_EXPAN0_reg_19_9_inst : FD1 port map( D => n5185, CP => CLK_I, Q => 
                           n_2844, QN => n2802);
   KEY_EXPAN0_reg_18_9_inst : FD1 port map( D => n5184, CP => CLK_I, Q => 
                           n_2845, QN => n2801);
   KEY_EXPAN0_reg_17_9_inst : FD1 port map( D => n5183, CP => CLK_I, Q => 
                           n_2846, QN => n2804);
   KEY_EXPAN0_reg_16_9_inst : FD1 port map( D => n5182, CP => CLK_I, Q => 
                           n_2847, QN => n2803);
   KEY_EXPAN0_reg_15_9_inst : FD1 port map( D => n5181, CP => CLK_I, Q => 
                           n_2848, QN => n2790);
   KEY_EXPAN0_reg_14_9_inst : FD1 port map( D => n5180, CP => CLK_I, Q => 
                           n_2849, QN => n2789);
   KEY_EXPAN0_reg_13_9_inst : FD1 port map( D => n5179, CP => CLK_I, Q => 
                           n_2850, QN => n2792);
   KEY_EXPAN0_reg_12_9_inst : FD1 port map( D => n5178, CP => CLK_I, Q => 
                           n_2851, QN => n2791);
   KEY_EXPAN0_reg_11_9_inst : FD1 port map( D => n5177, CP => CLK_I, Q => 
                           n_2852, QN => n2794);
   KEY_EXPAN0_reg_10_9_inst : FD1 port map( D => n5176, CP => CLK_I, Q => 
                           n_2853, QN => n2793);
   KEY_EXPAN0_reg_9_9_inst : FD1 port map( D => n5175, CP => CLK_I, Q => n_2854
                           , QN => n2796);
   KEY_EXPAN0_reg_8_9_inst : FD1 port map( D => n5174, CP => CLK_I, Q => n_2855
                           , QN => n2795);
   KEY_EXPAN0_reg_7_9_inst : FD1 port map( D => n5173, CP => CLK_I, Q => n_2856
                           , QN => n2782);
   KEY_EXPAN0_reg_6_9_inst : FD1 port map( D => n5172, CP => CLK_I, Q => n_2857
                           , QN => n2781);
   KEY_EXPAN0_reg_5_9_inst : FD1 port map( D => n5171, CP => CLK_I, Q => n_2858
                           , QN => n2784);
   KEY_EXPAN0_reg_4_9_inst : FD1 port map( D => n5170, CP => CLK_I, Q => n_2859
                           , QN => n2783);
   KEY_EXPAN0_reg_3_9_inst : FD1 port map( D => n5169, CP => CLK_I, Q => n_2860
                           , QN => n2786);
   KEY_EXPAN0_reg_2_9_inst : FD1 port map( D => n5168, CP => CLK_I, Q => n_2861
                           , QN => n2785);
   KEY_EXPAN0_reg_1_9_inst : FD1 port map( D => n5167, CP => CLK_I, Q => n_2862
                           , QN => n2788);
   KEY_EXPAN0_reg_0_9_inst : FD1 port map( D => n5166, CP => CLK_I, Q => n_2863
                           , QN => n2787);
   v_KEY_COL_OUT0_reg_9_inst : FD1 port map( D => n4553, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_9_port, QN => n1903);
   v_TEMP_VECTOR_reg_0_inst : FD1 port map( D => n6695, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_0_port, QN => n1992);
   KEY_EXPAN0_reg_63_0_inst : FD1 port map( D => n4653, CP => CLK_I, Q => 
                           n_2864, QN => n2709);
   KEY_EXPAN0_reg_62_0_inst : FD1 port map( D => n4652, CP => CLK_I, Q => 
                           n_2865, QN => n2708);
   KEY_EXPAN0_reg_61_0_inst : FD1 port map( D => n4651, CP => CLK_I, Q => 
                           n_2866, QN => n2711);
   KEY_EXPAN0_reg_60_0_inst : FD1 port map( D => n4650, CP => CLK_I, Q => 
                           n_2867, QN => n2710);
   KEY_EXPAN0_reg_59_0_inst : FD1 port map( D => n4649, CP => CLK_I, Q => 
                           n_2868, QN => n2713);
   KEY_EXPAN0_reg_58_0_inst : FD1 port map( D => n4648, CP => CLK_I, Q => 
                           n_2869, QN => n2712);
   KEY_EXPAN0_reg_57_0_inst : FD1 port map( D => n4647, CP => CLK_I, Q => 
                           n_2870, QN => n2715);
   KEY_EXPAN0_reg_56_0_inst : FD1 port map( D => n4646, CP => CLK_I, Q => 
                           n_2871, QN => n2714);
   KEY_EXPAN0_reg_55_0_inst : FD1 port map( D => n4645, CP => CLK_I, Q => 
                           n_2872, QN => n2701);
   KEY_EXPAN0_reg_54_0_inst : FD1 port map( D => n4644, CP => CLK_I, Q => 
                           n_2873, QN => n2700);
   KEY_EXPAN0_reg_53_0_inst : FD1 port map( D => n4643, CP => CLK_I, Q => 
                           n_2874, QN => n2703);
   KEY_EXPAN0_reg_52_0_inst : FD1 port map( D => n4642, CP => CLK_I, Q => 
                           n_2875, QN => n2702);
   KEY_EXPAN0_reg_51_0_inst : FD1 port map( D => n4641, CP => CLK_I, Q => 
                           n_2876, QN => n2705);
   KEY_EXPAN0_reg_50_0_inst : FD1 port map( D => n4640, CP => CLK_I, Q => 
                           n_2877, QN => n2704);
   KEY_EXPAN0_reg_49_0_inst : FD1 port map( D => n4639, CP => CLK_I, Q => 
                           n_2878, QN => n2707);
   KEY_EXPAN0_reg_48_0_inst : FD1 port map( D => n4638, CP => CLK_I, Q => 
                           n_2879, QN => n2706);
   KEY_EXPAN0_reg_47_0_inst : FD1 port map( D => n4637, CP => CLK_I, Q => 
                           n_2880, QN => n2693);
   KEY_EXPAN0_reg_46_0_inst : FD1 port map( D => n4636, CP => CLK_I, Q => 
                           n_2881, QN => n2692);
   KEY_EXPAN0_reg_45_0_inst : FD1 port map( D => n4635, CP => CLK_I, Q => 
                           n_2882, QN => n2695);
   KEY_EXPAN0_reg_44_0_inst : FD1 port map( D => n4634, CP => CLK_I, Q => 
                           n_2883, QN => n2694);
   KEY_EXPAN0_reg_43_0_inst : FD1 port map( D => n4633, CP => CLK_I, Q => 
                           n_2884, QN => n2697);
   KEY_EXPAN0_reg_42_0_inst : FD1 port map( D => n4632, CP => CLK_I, Q => 
                           n_2885, QN => n2696);
   KEY_EXPAN0_reg_41_0_inst : FD1 port map( D => n4631, CP => CLK_I, Q => 
                           n_2886, QN => n2699);
   KEY_EXPAN0_reg_40_0_inst : FD1 port map( D => n4630, CP => CLK_I, Q => 
                           n_2887, QN => n2698);
   KEY_EXPAN0_reg_39_0_inst : FD1 port map( D => n4629, CP => CLK_I, Q => 
                           n_2888, QN => n2685);
   KEY_EXPAN0_reg_38_0_inst : FD1 port map( D => n4628, CP => CLK_I, Q => 
                           n_2889, QN => n2684);
   KEY_EXPAN0_reg_37_0_inst : FD1 port map( D => n4627, CP => CLK_I, Q => 
                           n_2890, QN => n2687);
   KEY_EXPAN0_reg_36_0_inst : FD1 port map( D => n4626, CP => CLK_I, Q => 
                           n_2891, QN => n2686);
   KEY_EXPAN0_reg_35_0_inst : FD1 port map( D => n4625, CP => CLK_I, Q => 
                           n_2892, QN => n2689);
   KEY_EXPAN0_reg_34_0_inst : FD1 port map( D => n4624, CP => CLK_I, Q => 
                           n_2893, QN => n2688);
   KEY_EXPAN0_reg_33_0_inst : FD1 port map( D => n4623, CP => CLK_I, Q => 
                           n_2894, QN => n2691);
   KEY_EXPAN0_reg_32_0_inst : FD1 port map( D => n4622, CP => CLK_I, Q => 
                           n_2895, QN => n2690);
   KEY_EXPAN0_reg_31_0_inst : FD1 port map( D => n4621, CP => CLK_I, Q => 
                           n_2896, QN => n2741);
   KEY_EXPAN0_reg_30_0_inst : FD1 port map( D => n4620, CP => CLK_I, Q => 
                           n_2897, QN => n2740);
   KEY_EXPAN0_reg_29_0_inst : FD1 port map( D => n4619, CP => CLK_I, Q => 
                           n_2898, QN => n2743);
   KEY_EXPAN0_reg_28_0_inst : FD1 port map( D => n4618, CP => CLK_I, Q => 
                           n_2899, QN => n2742);
   KEY_EXPAN0_reg_27_0_inst : FD1 port map( D => n4617, CP => CLK_I, Q => 
                           n_2900, QN => n2745);
   KEY_EXPAN0_reg_26_0_inst : FD1 port map( D => n4616, CP => CLK_I, Q => 
                           n_2901, QN => n2744);
   KEY_EXPAN0_reg_25_0_inst : FD1 port map( D => n4615, CP => CLK_I, Q => 
                           n_2902, QN => n2747);
   KEY_EXPAN0_reg_24_0_inst : FD1 port map( D => n4614, CP => CLK_I, Q => 
                           n_2903, QN => n2746);
   KEY_EXPAN0_reg_23_0_inst : FD1 port map( D => n4613, CP => CLK_I, Q => 
                           n_2904, QN => n2733);
   KEY_EXPAN0_reg_22_0_inst : FD1 port map( D => n4612, CP => CLK_I, Q => 
                           n_2905, QN => n2732);
   KEY_EXPAN0_reg_21_0_inst : FD1 port map( D => n4611, CP => CLK_I, Q => 
                           n_2906, QN => n2735);
   KEY_EXPAN0_reg_20_0_inst : FD1 port map( D => n4610, CP => CLK_I, Q => 
                           n_2907, QN => n2734);
   KEY_EXPAN0_reg_19_0_inst : FD1 port map( D => n4609, CP => CLK_I, Q => 
                           n_2908, QN => n2737);
   KEY_EXPAN0_reg_18_0_inst : FD1 port map( D => n4608, CP => CLK_I, Q => 
                           n_2909, QN => n2736);
   KEY_EXPAN0_reg_17_0_inst : FD1 port map( D => n4607, CP => CLK_I, Q => 
                           n_2910, QN => n2739);
   KEY_EXPAN0_reg_16_0_inst : FD1 port map( D => n4606, CP => CLK_I, Q => 
                           n_2911, QN => n2738);
   KEY_EXPAN0_reg_15_0_inst : FD1 port map( D => n4605, CP => CLK_I, Q => 
                           n_2912, QN => n2725);
   KEY_EXPAN0_reg_14_0_inst : FD1 port map( D => n4604, CP => CLK_I, Q => 
                           n_2913, QN => n2724);
   KEY_EXPAN0_reg_13_0_inst : FD1 port map( D => n4603, CP => CLK_I, Q => 
                           n_2914, QN => n2727);
   KEY_EXPAN0_reg_12_0_inst : FD1 port map( D => n4602, CP => CLK_I, Q => 
                           n_2915, QN => n2726);
   KEY_EXPAN0_reg_11_0_inst : FD1 port map( D => n4601, CP => CLK_I, Q => 
                           n_2916, QN => n2729);
   KEY_EXPAN0_reg_10_0_inst : FD1 port map( D => n4600, CP => CLK_I, Q => 
                           n_2917, QN => n2728);
   KEY_EXPAN0_reg_9_0_inst : FD1 port map( D => n4599, CP => CLK_I, Q => n_2918
                           , QN => n2731);
   KEY_EXPAN0_reg_8_0_inst : FD1 port map( D => n4598, CP => CLK_I, Q => n_2919
                           , QN => n2730);
   KEY_EXPAN0_reg_7_0_inst : FD1 port map( D => n4597, CP => CLK_I, Q => n_2920
                           , QN => n2717);
   KEY_EXPAN0_reg_6_0_inst : FD1 port map( D => n4596, CP => CLK_I, Q => n_2921
                           , QN => n2716);
   KEY_EXPAN0_reg_5_0_inst : FD1 port map( D => n4595, CP => CLK_I, Q => n_2922
                           , QN => n2719);
   KEY_EXPAN0_reg_4_0_inst : FD1 port map( D => n4594, CP => CLK_I, Q => n_2923
                           , QN => n2718);
   KEY_EXPAN0_reg_3_0_inst : FD1 port map( D => n4593, CP => CLK_I, Q => n_2924
                           , QN => n2721);
   KEY_EXPAN0_reg_2_0_inst : FD1 port map( D => n4592, CP => CLK_I, Q => n_2925
                           , QN => n2720);
   KEY_EXPAN0_reg_1_0_inst : FD1 port map( D => n4591, CP => CLK_I, Q => n_2926
                           , QN => n2723);
   KEY_EXPAN0_reg_0_0_inst : FD1 port map( D => n4590, CP => CLK_I, Q => n_2927
                           , QN => n2722);
   v_KEY_COL_OUT0_reg_0_inst : FD1 port map( D => n4552, CP => CLK_I, Q => 
                           n2748, QN => n1887);
   v_TEMP_VECTOR_reg_24_inst : FD1 port map( D => n6671, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_24_port, QN => n_2928);
   KEY_EXPAN0_reg_63_24_inst : FD1 port map( D => n6189, CP => CLK_I, Q => 
                           n_2929, QN => n2645);
   KEY_EXPAN0_reg_62_24_inst : FD1 port map( D => n6188, CP => CLK_I, Q => 
                           n_2930, QN => n2644);
   KEY_EXPAN0_reg_61_24_inst : FD1 port map( D => n6187, CP => CLK_I, Q => 
                           n_2931, QN => n2647);
   KEY_EXPAN0_reg_60_24_inst : FD1 port map( D => n6186, CP => CLK_I, Q => 
                           n_2932, QN => n2646);
   KEY_EXPAN0_reg_59_24_inst : FD1 port map( D => n6185, CP => CLK_I, Q => 
                           n_2933, QN => n2649);
   KEY_EXPAN0_reg_58_24_inst : FD1 port map( D => n6184, CP => CLK_I, Q => 
                           n_2934, QN => n2648);
   KEY_EXPAN0_reg_57_24_inst : FD1 port map( D => n6183, CP => CLK_I, Q => 
                           n_2935, QN => n2651);
   KEY_EXPAN0_reg_56_24_inst : FD1 port map( D => n6182, CP => CLK_I, Q => 
                           n_2936, QN => n2650);
   KEY_EXPAN0_reg_55_24_inst : FD1 port map( D => n6181, CP => CLK_I, Q => 
                           n_2937, QN => n2637);
   KEY_EXPAN0_reg_54_24_inst : FD1 port map( D => n6180, CP => CLK_I, Q => 
                           n_2938, QN => n2636);
   KEY_EXPAN0_reg_53_24_inst : FD1 port map( D => n6179, CP => CLK_I, Q => 
                           n_2939, QN => n2639);
   KEY_EXPAN0_reg_52_24_inst : FD1 port map( D => n6178, CP => CLK_I, Q => 
                           n_2940, QN => n2638);
   KEY_EXPAN0_reg_51_24_inst : FD1 port map( D => n6177, CP => CLK_I, Q => 
                           n_2941, QN => n2641);
   KEY_EXPAN0_reg_50_24_inst : FD1 port map( D => n6176, CP => CLK_I, Q => 
                           n_2942, QN => n2640);
   KEY_EXPAN0_reg_49_24_inst : FD1 port map( D => n6175, CP => CLK_I, Q => 
                           n_2943, QN => n2643);
   KEY_EXPAN0_reg_48_24_inst : FD1 port map( D => n6174, CP => CLK_I, Q => 
                           n_2944, QN => n2642);
   KEY_EXPAN0_reg_47_24_inst : FD1 port map( D => n6173, CP => CLK_I, Q => 
                           n_2945, QN => n2629);
   KEY_EXPAN0_reg_46_24_inst : FD1 port map( D => n6172, CP => CLK_I, Q => 
                           n_2946, QN => n2628);
   KEY_EXPAN0_reg_45_24_inst : FD1 port map( D => n6171, CP => CLK_I, Q => 
                           n_2947, QN => n2631);
   KEY_EXPAN0_reg_44_24_inst : FD1 port map( D => n6170, CP => CLK_I, Q => 
                           n_2948, QN => n2630);
   KEY_EXPAN0_reg_43_24_inst : FD1 port map( D => n6169, CP => CLK_I, Q => 
                           n_2949, QN => n2633);
   KEY_EXPAN0_reg_42_24_inst : FD1 port map( D => n6168, CP => CLK_I, Q => 
                           n_2950, QN => n2632);
   KEY_EXPAN0_reg_41_24_inst : FD1 port map( D => n6167, CP => CLK_I, Q => 
                           n_2951, QN => n2635);
   KEY_EXPAN0_reg_40_24_inst : FD1 port map( D => n6166, CP => CLK_I, Q => 
                           n_2952, QN => n2634);
   KEY_EXPAN0_reg_39_24_inst : FD1 port map( D => n6165, CP => CLK_I, Q => 
                           n_2953, QN => n2621);
   KEY_EXPAN0_reg_38_24_inst : FD1 port map( D => n6164, CP => CLK_I, Q => 
                           n_2954, QN => n2620);
   KEY_EXPAN0_reg_37_24_inst : FD1 port map( D => n6163, CP => CLK_I, Q => 
                           n_2955, QN => n2623);
   KEY_EXPAN0_reg_36_24_inst : FD1 port map( D => n6162, CP => CLK_I, Q => 
                           n_2956, QN => n2622);
   KEY_EXPAN0_reg_35_24_inst : FD1 port map( D => n6161, CP => CLK_I, Q => 
                           n_2957, QN => n2625);
   KEY_EXPAN0_reg_34_24_inst : FD1 port map( D => n6160, CP => CLK_I, Q => 
                           n_2958, QN => n2624);
   KEY_EXPAN0_reg_33_24_inst : FD1 port map( D => n6159, CP => CLK_I, Q => 
                           n_2959, QN => n2627);
   KEY_EXPAN0_reg_32_24_inst : FD1 port map( D => n6158, CP => CLK_I, Q => 
                           n_2960, QN => n2626);
   KEY_EXPAN0_reg_31_24_inst : FD1 port map( D => n6157, CP => CLK_I, Q => 
                           n_2961, QN => n2677);
   KEY_EXPAN0_reg_30_24_inst : FD1 port map( D => n6156, CP => CLK_I, Q => 
                           n_2962, QN => n2676);
   KEY_EXPAN0_reg_29_24_inst : FD1 port map( D => n6155, CP => CLK_I, Q => 
                           n_2963, QN => n2679);
   KEY_EXPAN0_reg_28_24_inst : FD1 port map( D => n6154, CP => CLK_I, Q => 
                           n_2964, QN => n2678);
   KEY_EXPAN0_reg_27_24_inst : FD1 port map( D => n6153, CP => CLK_I, Q => 
                           n_2965, QN => n2681);
   KEY_EXPAN0_reg_26_24_inst : FD1 port map( D => n6152, CP => CLK_I, Q => 
                           n_2966, QN => n2680);
   KEY_EXPAN0_reg_25_24_inst : FD1 port map( D => n6151, CP => CLK_I, Q => 
                           n_2967, QN => n2683);
   KEY_EXPAN0_reg_24_24_inst : FD1 port map( D => n6150, CP => CLK_I, Q => 
                           n_2968, QN => n2682);
   KEY_EXPAN0_reg_23_24_inst : FD1 port map( D => n6149, CP => CLK_I, Q => 
                           n_2969, QN => n2669);
   KEY_EXPAN0_reg_22_24_inst : FD1 port map( D => n6148, CP => CLK_I, Q => 
                           n_2970, QN => n2668);
   KEY_EXPAN0_reg_21_24_inst : FD1 port map( D => n6147, CP => CLK_I, Q => 
                           n_2971, QN => n2671);
   KEY_EXPAN0_reg_20_24_inst : FD1 port map( D => n6146, CP => CLK_I, Q => 
                           n_2972, QN => n2670);
   KEY_EXPAN0_reg_19_24_inst : FD1 port map( D => n6145, CP => CLK_I, Q => 
                           n_2973, QN => n2673);
   KEY_EXPAN0_reg_18_24_inst : FD1 port map( D => n6144, CP => CLK_I, Q => 
                           n_2974, QN => n2672);
   KEY_EXPAN0_reg_17_24_inst : FD1 port map( D => n6143, CP => CLK_I, Q => 
                           n_2975, QN => n2675);
   KEY_EXPAN0_reg_16_24_inst : FD1 port map( D => n6142, CP => CLK_I, Q => 
                           n_2976, QN => n2674);
   KEY_EXPAN0_reg_15_24_inst : FD1 port map( D => n6141, CP => CLK_I, Q => 
                           n_2977, QN => n2661);
   KEY_EXPAN0_reg_14_24_inst : FD1 port map( D => n6140, CP => CLK_I, Q => 
                           n_2978, QN => n2660);
   KEY_EXPAN0_reg_13_24_inst : FD1 port map( D => n6139, CP => CLK_I, Q => 
                           n_2979, QN => n2663);
   KEY_EXPAN0_reg_12_24_inst : FD1 port map( D => n6138, CP => CLK_I, Q => 
                           n_2980, QN => n2662);
   KEY_EXPAN0_reg_11_24_inst : FD1 port map( D => n6137, CP => CLK_I, Q => 
                           n_2981, QN => n2665);
   KEY_EXPAN0_reg_10_24_inst : FD1 port map( D => n6136, CP => CLK_I, Q => 
                           n_2982, QN => n2664);
   KEY_EXPAN0_reg_9_24_inst : FD1 port map( D => n6135, CP => CLK_I, Q => 
                           n_2983, QN => n2667);
   KEY_EXPAN0_reg_8_24_inst : FD1 port map( D => n6134, CP => CLK_I, Q => 
                           n_2984, QN => n2666);
   KEY_EXPAN0_reg_7_24_inst : FD1 port map( D => n6133, CP => CLK_I, Q => 
                           n_2985, QN => n2653);
   KEY_EXPAN0_reg_6_24_inst : FD1 port map( D => n6132, CP => CLK_I, Q => 
                           n_2986, QN => n2652);
   KEY_EXPAN0_reg_5_24_inst : FD1 port map( D => n6131, CP => CLK_I, Q => 
                           n_2987, QN => n2655);
   KEY_EXPAN0_reg_4_24_inst : FD1 port map( D => n6130, CP => CLK_I, Q => 
                           n_2988, QN => n2654);
   KEY_EXPAN0_reg_3_24_inst : FD1 port map( D => n6129, CP => CLK_I, Q => 
                           n_2989, QN => n2657);
   KEY_EXPAN0_reg_2_24_inst : FD1 port map( D => n6128, CP => CLK_I, Q => 
                           n_2990, QN => n2656);
   KEY_EXPAN0_reg_1_24_inst : FD1 port map( D => n6127, CP => CLK_I, Q => 
                           n_2991, QN => n2659);
   KEY_EXPAN0_reg_0_24_inst : FD1 port map( D => n6126, CP => CLK_I, Q => 
                           n_2992, QN => n2658);
   v_KEY_COL_OUT0_reg_24_inst : FD1 port map( D => n4551, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_24_port, QN => n355);
   v_TEMP_VECTOR_reg_16_inst : FD1 port map( D => n6679, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_16_port, QN => n_2993);
   KEY_EXPAN0_reg_63_16_inst : FD1 port map( D => n5677, CP => CLK_I, Q => 
                           n_2994, QN => n2581);
   KEY_EXPAN0_reg_62_16_inst : FD1 port map( D => n5676, CP => CLK_I, Q => 
                           n_2995, QN => n2580);
   KEY_EXPAN0_reg_61_16_inst : FD1 port map( D => n5675, CP => CLK_I, Q => 
                           n_2996, QN => n2583);
   KEY_EXPAN0_reg_60_16_inst : FD1 port map( D => n5674, CP => CLK_I, Q => 
                           n_2997, QN => n2582);
   KEY_EXPAN0_reg_59_16_inst : FD1 port map( D => n5673, CP => CLK_I, Q => 
                           n_2998, QN => n2585);
   KEY_EXPAN0_reg_58_16_inst : FD1 port map( D => n5672, CP => CLK_I, Q => 
                           n_2999, QN => n2584);
   KEY_EXPAN0_reg_57_16_inst : FD1 port map( D => n5671, CP => CLK_I, Q => 
                           n_3000, QN => n2587);
   KEY_EXPAN0_reg_56_16_inst : FD1 port map( D => n5670, CP => CLK_I, Q => 
                           n_3001, QN => n2586);
   KEY_EXPAN0_reg_55_16_inst : FD1 port map( D => n5669, CP => CLK_I, Q => 
                           n_3002, QN => n2573);
   KEY_EXPAN0_reg_54_16_inst : FD1 port map( D => n5668, CP => CLK_I, Q => 
                           n_3003, QN => n2572);
   KEY_EXPAN0_reg_53_16_inst : FD1 port map( D => n5667, CP => CLK_I, Q => 
                           n_3004, QN => n2575);
   KEY_EXPAN0_reg_52_16_inst : FD1 port map( D => n5666, CP => CLK_I, Q => 
                           n_3005, QN => n2574);
   KEY_EXPAN0_reg_51_16_inst : FD1 port map( D => n5665, CP => CLK_I, Q => 
                           n_3006, QN => n2577);
   KEY_EXPAN0_reg_50_16_inst : FD1 port map( D => n5664, CP => CLK_I, Q => 
                           n_3007, QN => n2576);
   KEY_EXPAN0_reg_49_16_inst : FD1 port map( D => n5663, CP => CLK_I, Q => 
                           n_3008, QN => n2579);
   KEY_EXPAN0_reg_48_16_inst : FD1 port map( D => n5662, CP => CLK_I, Q => 
                           n_3009, QN => n2578);
   KEY_EXPAN0_reg_47_16_inst : FD1 port map( D => n5661, CP => CLK_I, Q => 
                           n_3010, QN => n2565);
   KEY_EXPAN0_reg_46_16_inst : FD1 port map( D => n5660, CP => CLK_I, Q => 
                           n_3011, QN => n2564);
   KEY_EXPAN0_reg_45_16_inst : FD1 port map( D => n5659, CP => CLK_I, Q => 
                           n_3012, QN => n2567);
   KEY_EXPAN0_reg_44_16_inst : FD1 port map( D => n5658, CP => CLK_I, Q => 
                           n_3013, QN => n2566);
   KEY_EXPAN0_reg_43_16_inst : FD1 port map( D => n5657, CP => CLK_I, Q => 
                           n_3014, QN => n2569);
   KEY_EXPAN0_reg_42_16_inst : FD1 port map( D => n5656, CP => CLK_I, Q => 
                           n_3015, QN => n2568);
   KEY_EXPAN0_reg_41_16_inst : FD1 port map( D => n5655, CP => CLK_I, Q => 
                           n_3016, QN => n2571);
   KEY_EXPAN0_reg_40_16_inst : FD1 port map( D => n5654, CP => CLK_I, Q => 
                           n_3017, QN => n2570);
   KEY_EXPAN0_reg_39_16_inst : FD1 port map( D => n5653, CP => CLK_I, Q => 
                           n_3018, QN => n2557);
   KEY_EXPAN0_reg_38_16_inst : FD1 port map( D => n5652, CP => CLK_I, Q => 
                           n_3019, QN => n2556);
   KEY_EXPAN0_reg_37_16_inst : FD1 port map( D => n5651, CP => CLK_I, Q => 
                           n_3020, QN => n2559);
   KEY_EXPAN0_reg_36_16_inst : FD1 port map( D => n5650, CP => CLK_I, Q => 
                           n_3021, QN => n2558);
   KEY_EXPAN0_reg_35_16_inst : FD1 port map( D => n5649, CP => CLK_I, Q => 
                           n_3022, QN => n2561);
   KEY_EXPAN0_reg_34_16_inst : FD1 port map( D => n5648, CP => CLK_I, Q => 
                           n_3023, QN => n2560);
   KEY_EXPAN0_reg_33_16_inst : FD1 port map( D => n5647, CP => CLK_I, Q => 
                           n_3024, QN => n2563);
   KEY_EXPAN0_reg_32_16_inst : FD1 port map( D => n5646, CP => CLK_I, Q => 
                           n_3025, QN => n2562);
   KEY_EXPAN0_reg_31_16_inst : FD1 port map( D => n5645, CP => CLK_I, Q => 
                           n_3026, QN => n2613);
   KEY_EXPAN0_reg_30_16_inst : FD1 port map( D => n5644, CP => CLK_I, Q => 
                           n_3027, QN => n2612);
   KEY_EXPAN0_reg_29_16_inst : FD1 port map( D => n5643, CP => CLK_I, Q => 
                           n_3028, QN => n2615);
   KEY_EXPAN0_reg_28_16_inst : FD1 port map( D => n5642, CP => CLK_I, Q => 
                           n_3029, QN => n2614);
   KEY_EXPAN0_reg_27_16_inst : FD1 port map( D => n5641, CP => CLK_I, Q => 
                           n_3030, QN => n2617);
   KEY_EXPAN0_reg_26_16_inst : FD1 port map( D => n5640, CP => CLK_I, Q => 
                           n_3031, QN => n2616);
   KEY_EXPAN0_reg_25_16_inst : FD1 port map( D => n5639, CP => CLK_I, Q => 
                           n_3032, QN => n2619);
   KEY_EXPAN0_reg_24_16_inst : FD1 port map( D => n5638, CP => CLK_I, Q => 
                           n_3033, QN => n2618);
   KEY_EXPAN0_reg_23_16_inst : FD1 port map( D => n5637, CP => CLK_I, Q => 
                           n_3034, QN => n2605);
   KEY_EXPAN0_reg_22_16_inst : FD1 port map( D => n5636, CP => CLK_I, Q => 
                           n_3035, QN => n2604);
   KEY_EXPAN0_reg_21_16_inst : FD1 port map( D => n5635, CP => CLK_I, Q => 
                           n_3036, QN => n2607);
   KEY_EXPAN0_reg_20_16_inst : FD1 port map( D => n5634, CP => CLK_I, Q => 
                           n_3037, QN => n2606);
   KEY_EXPAN0_reg_19_16_inst : FD1 port map( D => n5633, CP => CLK_I, Q => 
                           n_3038, QN => n2609);
   KEY_EXPAN0_reg_18_16_inst : FD1 port map( D => n5632, CP => CLK_I, Q => 
                           n_3039, QN => n2608);
   KEY_EXPAN0_reg_17_16_inst : FD1 port map( D => n5631, CP => CLK_I, Q => 
                           n_3040, QN => n2611);
   KEY_EXPAN0_reg_16_16_inst : FD1 port map( D => n5630, CP => CLK_I, Q => 
                           n_3041, QN => n2610);
   KEY_EXPAN0_reg_15_16_inst : FD1 port map( D => n5629, CP => CLK_I, Q => 
                           n_3042, QN => n2597);
   KEY_EXPAN0_reg_14_16_inst : FD1 port map( D => n5628, CP => CLK_I, Q => 
                           n_3043, QN => n2596);
   KEY_EXPAN0_reg_13_16_inst : FD1 port map( D => n5627, CP => CLK_I, Q => 
                           n_3044, QN => n2599);
   KEY_EXPAN0_reg_12_16_inst : FD1 port map( D => n5626, CP => CLK_I, Q => 
                           n_3045, QN => n2598);
   KEY_EXPAN0_reg_11_16_inst : FD1 port map( D => n5625, CP => CLK_I, Q => 
                           n_3046, QN => n2601);
   KEY_EXPAN0_reg_10_16_inst : FD1 port map( D => n5624, CP => CLK_I, Q => 
                           n_3047, QN => n2600);
   KEY_EXPAN0_reg_9_16_inst : FD1 port map( D => n5623, CP => CLK_I, Q => 
                           n_3048, QN => n2603);
   KEY_EXPAN0_reg_8_16_inst : FD1 port map( D => n5622, CP => CLK_I, Q => 
                           n_3049, QN => n2602);
   KEY_EXPAN0_reg_7_16_inst : FD1 port map( D => n5621, CP => CLK_I, Q => 
                           n_3050, QN => n2589);
   KEY_EXPAN0_reg_6_16_inst : FD1 port map( D => n5620, CP => CLK_I, Q => 
                           n_3051, QN => n2588);
   KEY_EXPAN0_reg_5_16_inst : FD1 port map( D => n5619, CP => CLK_I, Q => 
                           n_3052, QN => n2591);
   KEY_EXPAN0_reg_4_16_inst : FD1 port map( D => n5618, CP => CLK_I, Q => 
                           n_3053, QN => n2590);
   KEY_EXPAN0_reg_3_16_inst : FD1 port map( D => n5617, CP => CLK_I, Q => 
                           n_3054, QN => n2593);
   KEY_EXPAN0_reg_2_16_inst : FD1 port map( D => n5616, CP => CLK_I, Q => 
                           n_3055, QN => n2592);
   KEY_EXPAN0_reg_1_16_inst : FD1 port map( D => n5615, CP => CLK_I, Q => 
                           n_3056, QN => n2595);
   KEY_EXPAN0_reg_0_16_inst : FD1 port map( D => n5614, CP => CLK_I, Q => 
                           n_3057, QN => n2594);
   v_KEY_COL_OUT0_reg_16_inst : FD1 port map( D => n4550, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_16_port, QN => n388);
   v_TEMP_VECTOR_reg_8_inst : FD1 port map( D => n6687, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_8_port, QN => n_3058);
   KEY_EXPAN0_reg_63_8_inst : FD1 port map( D => n5165, CP => CLK_I, Q => 
                           n_3059, QN => n2517);
   KEY_EXPAN0_reg_62_8_inst : FD1 port map( D => n5164, CP => CLK_I, Q => 
                           n_3060, QN => n2516);
   KEY_EXPAN0_reg_61_8_inst : FD1 port map( D => n5163, CP => CLK_I, Q => 
                           n_3061, QN => n2519);
   KEY_EXPAN0_reg_60_8_inst : FD1 port map( D => n5162, CP => CLK_I, Q => 
                           n_3062, QN => n2518);
   KEY_EXPAN0_reg_59_8_inst : FD1 port map( D => n5161, CP => CLK_I, Q => 
                           n_3063, QN => n2521);
   KEY_EXPAN0_reg_58_8_inst : FD1 port map( D => n5160, CP => CLK_I, Q => 
                           n_3064, QN => n2520);
   KEY_EXPAN0_reg_57_8_inst : FD1 port map( D => n5159, CP => CLK_I, Q => 
                           n_3065, QN => n2523);
   KEY_EXPAN0_reg_56_8_inst : FD1 port map( D => n5158, CP => CLK_I, Q => 
                           n_3066, QN => n2522);
   KEY_EXPAN0_reg_55_8_inst : FD1 port map( D => n5157, CP => CLK_I, Q => 
                           n_3067, QN => n2509);
   KEY_EXPAN0_reg_54_8_inst : FD1 port map( D => n5156, CP => CLK_I, Q => 
                           n_3068, QN => n2508);
   KEY_EXPAN0_reg_53_8_inst : FD1 port map( D => n5155, CP => CLK_I, Q => 
                           n_3069, QN => n2511);
   KEY_EXPAN0_reg_52_8_inst : FD1 port map( D => n5154, CP => CLK_I, Q => 
                           n_3070, QN => n2510);
   KEY_EXPAN0_reg_51_8_inst : FD1 port map( D => n5153, CP => CLK_I, Q => 
                           n_3071, QN => n2513);
   KEY_EXPAN0_reg_50_8_inst : FD1 port map( D => n5152, CP => CLK_I, Q => 
                           n_3072, QN => n2512);
   KEY_EXPAN0_reg_49_8_inst : FD1 port map( D => n5151, CP => CLK_I, Q => 
                           n_3073, QN => n2515);
   KEY_EXPAN0_reg_48_8_inst : FD1 port map( D => n5150, CP => CLK_I, Q => 
                           n_3074, QN => n2514);
   KEY_EXPAN0_reg_47_8_inst : FD1 port map( D => n5149, CP => CLK_I, Q => 
                           n_3075, QN => n2501);
   KEY_EXPAN0_reg_46_8_inst : FD1 port map( D => n5148, CP => CLK_I, Q => 
                           n_3076, QN => n2500);
   KEY_EXPAN0_reg_45_8_inst : FD1 port map( D => n5147, CP => CLK_I, Q => 
                           n_3077, QN => n2503);
   KEY_EXPAN0_reg_44_8_inst : FD1 port map( D => n5146, CP => CLK_I, Q => 
                           n_3078, QN => n2502);
   KEY_EXPAN0_reg_43_8_inst : FD1 port map( D => n5145, CP => CLK_I, Q => 
                           n_3079, QN => n2505);
   KEY_EXPAN0_reg_42_8_inst : FD1 port map( D => n5144, CP => CLK_I, Q => 
                           n_3080, QN => n2504);
   KEY_EXPAN0_reg_41_8_inst : FD1 port map( D => n5143, CP => CLK_I, Q => 
                           n_3081, QN => n2507);
   KEY_EXPAN0_reg_40_8_inst : FD1 port map( D => n5142, CP => CLK_I, Q => 
                           n_3082, QN => n2506);
   KEY_EXPAN0_reg_39_8_inst : FD1 port map( D => n5141, CP => CLK_I, Q => 
                           n_3083, QN => n2493);
   KEY_EXPAN0_reg_38_8_inst : FD1 port map( D => n5140, CP => CLK_I, Q => 
                           n_3084, QN => n2492);
   KEY_EXPAN0_reg_37_8_inst : FD1 port map( D => n5139, CP => CLK_I, Q => 
                           n_3085, QN => n2495);
   KEY_EXPAN0_reg_36_8_inst : FD1 port map( D => n5138, CP => CLK_I, Q => 
                           n_3086, QN => n2494);
   KEY_EXPAN0_reg_35_8_inst : FD1 port map( D => n5137, CP => CLK_I, Q => 
                           n_3087, QN => n2497);
   KEY_EXPAN0_reg_34_8_inst : FD1 port map( D => n5136, CP => CLK_I, Q => 
                           n_3088, QN => n2496);
   KEY_EXPAN0_reg_33_8_inst : FD1 port map( D => n5135, CP => CLK_I, Q => 
                           n_3089, QN => n2499);
   KEY_EXPAN0_reg_32_8_inst : FD1 port map( D => n5134, CP => CLK_I, Q => 
                           n_3090, QN => n2498);
   KEY_EXPAN0_reg_31_8_inst : FD1 port map( D => n5133, CP => CLK_I, Q => 
                           n_3091, QN => n2549);
   KEY_EXPAN0_reg_30_8_inst : FD1 port map( D => n5132, CP => CLK_I, Q => 
                           n_3092, QN => n2548);
   KEY_EXPAN0_reg_29_8_inst : FD1 port map( D => n5131, CP => CLK_I, Q => 
                           n_3093, QN => n2551);
   KEY_EXPAN0_reg_28_8_inst : FD1 port map( D => n5130, CP => CLK_I, Q => 
                           n_3094, QN => n2550);
   KEY_EXPAN0_reg_27_8_inst : FD1 port map( D => n5129, CP => CLK_I, Q => 
                           n_3095, QN => n2553);
   KEY_EXPAN0_reg_26_8_inst : FD1 port map( D => n5128, CP => CLK_I, Q => 
                           n_3096, QN => n2552);
   KEY_EXPAN0_reg_25_8_inst : FD1 port map( D => n5127, CP => CLK_I, Q => 
                           n_3097, QN => n2555);
   KEY_EXPAN0_reg_24_8_inst : FD1 port map( D => n5126, CP => CLK_I, Q => 
                           n_3098, QN => n2554);
   KEY_EXPAN0_reg_23_8_inst : FD1 port map( D => n5125, CP => CLK_I, Q => 
                           n_3099, QN => n2541);
   KEY_EXPAN0_reg_22_8_inst : FD1 port map( D => n5124, CP => CLK_I, Q => 
                           n_3100, QN => n2540);
   KEY_EXPAN0_reg_21_8_inst : FD1 port map( D => n5123, CP => CLK_I, Q => 
                           n_3101, QN => n2543);
   KEY_EXPAN0_reg_20_8_inst : FD1 port map( D => n5122, CP => CLK_I, Q => 
                           n_3102, QN => n2542);
   KEY_EXPAN0_reg_19_8_inst : FD1 port map( D => n5121, CP => CLK_I, Q => 
                           n_3103, QN => n2545);
   KEY_EXPAN0_reg_18_8_inst : FD1 port map( D => n5120, CP => CLK_I, Q => 
                           n_3104, QN => n2544);
   KEY_EXPAN0_reg_17_8_inst : FD1 port map( D => n5119, CP => CLK_I, Q => 
                           n_3105, QN => n2547);
   KEY_EXPAN0_reg_16_8_inst : FD1 port map( D => n5118, CP => CLK_I, Q => 
                           n_3106, QN => n2546);
   KEY_EXPAN0_reg_15_8_inst : FD1 port map( D => n5117, CP => CLK_I, Q => 
                           n_3107, QN => n2533);
   KEY_EXPAN0_reg_14_8_inst : FD1 port map( D => n5116, CP => CLK_I, Q => 
                           n_3108, QN => n2532);
   KEY_EXPAN0_reg_13_8_inst : FD1 port map( D => n5115, CP => CLK_I, Q => 
                           n_3109, QN => n2535);
   KEY_EXPAN0_reg_12_8_inst : FD1 port map( D => n5114, CP => CLK_I, Q => 
                           n_3110, QN => n2534);
   KEY_EXPAN0_reg_11_8_inst : FD1 port map( D => n5113, CP => CLK_I, Q => 
                           n_3111, QN => n2537);
   KEY_EXPAN0_reg_10_8_inst : FD1 port map( D => n5112, CP => CLK_I, Q => 
                           n_3112, QN => n2536);
   KEY_EXPAN0_reg_9_8_inst : FD1 port map( D => n5111, CP => CLK_I, Q => n_3113
                           , QN => n2539);
   KEY_EXPAN0_reg_8_8_inst : FD1 port map( D => n5110, CP => CLK_I, Q => n_3114
                           , QN => n2538);
   KEY_EXPAN0_reg_7_8_inst : FD1 port map( D => n5109, CP => CLK_I, Q => n_3115
                           , QN => n2525);
   KEY_EXPAN0_reg_6_8_inst : FD1 port map( D => n5108, CP => CLK_I, Q => n_3116
                           , QN => n2524);
   KEY_EXPAN0_reg_5_8_inst : FD1 port map( D => n5107, CP => CLK_I, Q => n_3117
                           , QN => n2527);
   KEY_EXPAN0_reg_4_8_inst : FD1 port map( D => n5106, CP => CLK_I, Q => n_3118
                           , QN => n2526);
   KEY_EXPAN0_reg_3_8_inst : FD1 port map( D => n5105, CP => CLK_I, Q => n_3119
                           , QN => n2529);
   KEY_EXPAN0_reg_2_8_inst : FD1 port map( D => n5104, CP => CLK_I, Q => n_3120
                           , QN => n2528);
   KEY_EXPAN0_reg_1_8_inst : FD1 port map( D => n5103, CP => CLK_I, Q => n_3121
                           , QN => n2531);
   KEY_EXPAN0_reg_0_8_inst : FD1 port map( D => n5102, CP => CLK_I, Q => n_3122
                           , QN => n2530);
   v_KEY_COL_OUT0_reg_8_inst : FD1 port map( D => n4549, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_8_port, QN => n394);
   U149 : OR3 port map( A => n155, B => n156, C => n157, Z => n66);
   U206 : OR3 port map( A => n6663, B => n363, C => n1918, Z => n223);
   U211 : OR2 port map( A => n6659, B => RESET_I, Z => n56);
   U215 : AN3 port map( A => n6662, B => n6663, C => n6661, Z => n230);
   U282 : AN3 port map( A => n363, B => n290, C => n6661, Z => n207);
   U293 : AN3 port map( A => n1918, B => n363, C => n290, Z => n280);
   U1923 : OR3 port map( A => n1878, B => n1929, C => n1930, Z => n1891);
   U2063 : AN3 port map( A => n1934, B => n1973, C => n267, Z => n2148);
   U2102 : OR3 port map( A => n377, B => n8247, C => n1951, Z => n2171);
   U2146 : AN3 port map( A => n2205, B => n1941, C => n2029, Z => n2194);
   U2165 : AN3 port map( A => n2082, B => n2147, C => n267, Z => n2217);
   U2166 : AN3 port map( A => n8263, B => n1957, C => n377, Z => n2216);
   U2209 : OR3 port map( A => n2072, B => n2206, C => n2174, Z => n2080);
   U2347 : AN3 port map( A => n2283, B => n366, C => n8282, Z => n175);
   U4494 : AN3 port map( A => n6639, B => n6640, C => n2469, Z => n2468);
   U4519 : AN3 port map( A => n6639, B => i_SRAM_ADDR_WR0_3_port, C => n2469, Z
                           => n2470);
   U4544 : AN3 port map( A => n6640, B => i_SRAM_ADDR_WR0_4_port, C => n2469, Z
                           => n2471);
   U4548 : AN3 port map( A => n6642, B => n6643, C => n6641, Z => n2452);
   U4552 : AN3 port map( A => n6642, B => i_SRAM_ADDR_WR0_0_port, C => n6641, Z
                           => n2454);
   U4556 : AN3 port map( A => n6643, B => i_SRAM_ADDR_WR0_1_port, C => n6641, Z
                           => n2455);
   U4560 : AN3 port map( A => i_SRAM_ADDR_WR0_0_port, B => 
                           i_SRAM_ADDR_WR0_1_port, C => n6641, Z => n2456);
   U4578 : AN4 port map( A => n2285, B => n2476, C => n2477, D => n2478, Z => 
                           n2475);
   U4582 : OR3 port map( A => n8280, B => n2305, C => n2111, Z => n2477);
   U4594 : AN3 port map( A => i_SRAM_ADDR_WR0_3_port, B => 
                           i_SRAM_ADDR_WR0_4_port, C => n2469, Z => n2472);
   U7 : NR2I port map( A => v_TEMP_VECTOR_31_port, B => n2304, Z => n19);
   U12 : NR2I port map( A => v_TEMP_VECTOR_30_port, B => n2304, Z => n26);
   U17 : NR2I port map( A => v_TEMP_VECTOR_29_port, B => n2304, Z => n31);
   U22 : NR2I port map( A => v_TEMP_VECTOR_28_port, B => n2304, Z => n36);
   U27 : NR2I port map( A => v_TEMP_VECTOR_27_port, B => n2304, Z => n41);
   U32 : NR2I port map( A => v_TEMP_VECTOR_26_port, B => n2304, Z => n46);
   U37 : NR2I port map( A => v_TEMP_VECTOR_25_port, B => n2304, Z => n51);
   U40 : NR2I port map( A => n56, B => n57, Z => n18);
   U41 : NR2I port map( A => n58, B => n8221, Z => n17);
   U45 : NR2I port map( A => v_TEMP_VECTOR_24_port, B => n2304, Z => n60);
   U48 : ND2I port map( A => n64, B => n62, Z => n13);
   U49 : NR2I port map( A => n57, B => n65, Z => n64);
   U52 : ND2I port map( A => n8289, B => n1985, Z => n70);
   U57 : NR2I port map( A => v_TEMP_VECTOR_23_port, B => n2302, Z => n78);
   U62 : NR2I port map( A => v_TEMP_VECTOR_22_port, B => n2302, Z => n84);
   U67 : NR2I port map( A => v_TEMP_VECTOR_21_port, B => n2302, Z => n88);
   U72 : NR2I port map( A => v_TEMP_VECTOR_20_port, B => n2302, Z => n92);
   U77 : NR2I port map( A => v_TEMP_VECTOR_19_port, B => n2302, Z => n96);
   U82 : NR2I port map( A => v_TEMP_VECTOR_18_port, B => n2302, Z => n100);
   U87 : NR2I port map( A => v_TEMP_VECTOR_17_port, B => n2302, Z => n104);
   U90 : NR2I port map( A => n108, B => n56, Z => n77);
   U91 : NR2I port map( A => n8278, B => n58, Z => n76);
   U95 : NR2I port map( A => v_TEMP_VECTOR_16_port, B => n2302, Z => n110);
   U98 : ND2I port map( A => n113, B => n2166, Z => n73);
   U99 : NR2I port map( A => n108, B => n65, Z => n113);
   U105 : NR2I port map( A => v_TEMP_VECTOR_15_port, B => n2300, Z => n119);
   U110 : NR2I port map( A => v_TEMP_VECTOR_14_port, B => n2300, Z => n125);
   U115 : NR2I port map( A => v_TEMP_VECTOR_13_port, B => n2300, Z => n129);
   U120 : NR2I port map( A => v_TEMP_VECTOR_12_port, B => n2300, Z => n133);
   U125 : NR2I port map( A => v_TEMP_VECTOR_11_port, B => n2300, Z => n137);
   U130 : NR2I port map( A => v_TEMP_VECTOR_10_port, B => n2300, Z => n141);
   U135 : NR2I port map( A => v_TEMP_VECTOR_9_port, B => n2300, Z => n145);
   U138 : NR2I port map( A => n149, B => n56, Z => n118);
   U139 : NR2I port map( A => n8276, B => n58, Z => n117);
   U143 : NR2I port map( A => v_TEMP_VECTOR_8_port, B => n2300, Z => n151);
   U146 : ND2I port map( A => n154, B => n2168, Z => n114);
   U147 : NR2I port map( A => n149, B => n65, Z => n154);
   U152 : ND2I port map( A => n2297, B => n165, Z => n160);
   U154 : EOI port map( A => v_TEMP_VECTOR_7_port, B => n354, Z => n167);
   U156 : EOI port map( A => v_TEMP_VECTOR_15_port, B => n8287, Z => n158);
   U161 : ENI port map( A => n180, B => v_TEMP_VECTOR_14_port, Z => n179);
   U163 : EOI port map( A => v_TEMP_VECTOR_6_port, B => n4285, Z => n178);
   U167 : ND2I port map( A => n2297, B => n186, Z => n184);
   U169 : EOI port map( A => v_TEMP_VECTOR_5_port, B => n382, Z => n187);
   U171 : ENI port map( A => v_TEMP_VECTOR_13_port, B => n189, Z => n183);
   U175 : ND2I port map( A => n2297, B => n194, Z => n192);
   U177 : EOI port map( A => v_TEMP_VECTOR_4_port, B => n1630, Z => n195);
   U179 : ENI port map( A => n197, B => v_TEMP_VECTOR_12_port, Z => n191);
   U183 : ND2I port map( A => n2297, B => n202, Z => n200);
   U185 : EOI port map( A => v_TEMP_VECTOR_3_port, B => n1586, Z => n203);
   U187 : EOI port map( A => n205, B => v_TEMP_VECTOR_11_port, Z => n199);
   U191 : ND2I port map( A => n2297, B => n211, Z => n209);
   U193 : EOI port map( A => v_TEMP_VECTOR_2_port, B => n403, Z => n212);
   U195 : ENI port map( A => n214, B => v_TEMP_VECTOR_10_port, Z => n208);
   U197 : ND2I port map( A => n6661, B => n363, Z => n215);
   U200 : ND2I port map( A => n2297, B => n219, Z => n217);
   U202 : ND2I port map( A => n2140, B => n58, Z => n168);
   U203 : EOI port map( A => v_TEMP_VECTOR_1_port, B => n1542, Z => n220);
   U204 : ENI port map( A => n222, B => v_TEMP_VECTOR_9_port, Z => n216);
   U205 : ND2I port map( A => n6660, B => n223, Z => n222);
   U207 : ND2I port map( A => n2297, B => n8281, Z => n159);
   U210 : NR2I port map( A => n56, B => n8279, Z => n162);
   U214 : EOI port map( A => v_TEMP_VECTOR_8_port, B => n230, Z => n229);
   U216 : EOI port map( A => v_TEMP_VECTOR_0_port, B => n2748, Z => n228);
   U217 : NR2I port map( A => n8281, B => n231, Z => n177);
   U218 : NR2I port map( A => n65, B => n8279, Z => n164);
   U235 : ND2I port map( A => n245, B => n237, Z => n239);
   U237 : ND2I port map( A => n246, B => n8297, Z => n237);
   U241 : ND2I port map( A => n358, B => n288, Z => n253);
   U244 : ND2I port map( A => n259, B => n366, Z => n258);
   U256 : ND2I port map( A => n245, B => n260, Z => n262);
   U263 : ND2I port map( A => n8282, B => n8289, Z => n58);
   U266 : ND2I port map( A => n272, B => n8300, Z => n275);
   U268 : ND2I port map( A => n8215, B => n8300, Z => n277);
   U270 : ND2I port map( A => n278, B => n279, Z => n272);
   U273 : ND2I port map( A => n281, B => n8300, Z => n282);
   U275 : ND2I port map( A => n278, B => n284, Z => n281);
   U279 : NR2I port map( A => n4548, B => VALID_KEY_I, Z => n283);
   U283 : ND2I port map( A => n6662, B => n1918, Z => n190);
   U286 : ND2I port map( A => n6662, B => n290, Z => n289);
   U292 : ND2I port map( A => n6660, B => n280, Z => n291);
   U298 : NR2I port map( A => n293, B => n65, Z => n286);
   U300 : ND2I port map( A => n8286, B => n8164, Z => n67);
   U338 : ND2I port map( A => n315, B => n2488, Z => n307);
   U356 : ND2I port map( A => n315, B => n2487, Z => n318);
   U377 : ND2I port map( A => n8299, B => n288, Z => n338);
   U382 : NR2I port map( A => n341, B => n342, Z => n340);
   U426 : NR2I port map( A => n449, B => n450, Z => n448);
   U470 : NR2I port map( A => n493, B => n494, Z => n492);
   U514 : NR2I port map( A => n537, B => n538, Z => n536);
   U558 : NR2I port map( A => n581, B => n582, Z => n580);
   U602 : NR2I port map( A => n625, B => n626, Z => n624);
   U646 : NR2I port map( A => n669, B => n670, Z => n668);
   U690 : NR2I port map( A => n712, B => n713, Z => n711);
   U734 : NR2I port map( A => n756, B => n757, Z => n755);
   U778 : NR2I port map( A => n800, B => n801, Z => n799);
   U822 : NR2I port map( A => n844, B => n845, Z => n843);
   U866 : NR2I port map( A => n887, B => n888, Z => n886);
   U910 : NR2I port map( A => n931, B => n932, Z => n930);
   U954 : NR2I port map( A => n975, B => n976, Z => n974);
   U998 : NR2I port map( A => n1019, B => n1020, Z => n1018);
   U1042 : NR2I port map( A => n1062, B => n1063, Z => n1061);
   U1086 : NR2I port map( A => n1106, B => n1107, Z => n1105);
   U1130 : NR2I port map( A => n1150, B => n1151, Z => n1149);
   U1174 : NR2I port map( A => n1194, B => n1195, Z => n1193);
   U1218 : NR2I port map( A => n1237, B => n1238, Z => n1236);
   U1262 : NR2I port map( A => n1281, B => n1282, Z => n1280);
   U1306 : NR2I port map( A => n1325, B => n1326, Z => n1324);
   U1350 : NR2I port map( A => n1369, B => n1370, Z => n1368);
   U1394 : NR2I port map( A => n1412, B => n1413, Z => n1411);
   U1438 : NR2I port map( A => n1456, B => n1457, Z => n1455);
   U1482 : NR2I port map( A => n1500, B => n1501, Z => n1499);
   U1526 : NR2I port map( A => n1544, B => n1545, Z => n1543);
   U1570 : NR2I port map( A => n1588, B => n1589, Z => n1587);
   U1614 : NR2I port map( A => n1632, B => n1633, Z => n1631);
   U1658 : NR2I port map( A => n1676, B => n1677, Z => n1675);
   U1702 : NR2I port map( A => n1720, B => n1721, Z => n1719);
   U1746 : NR2I port map( A => n1763, B => n1764, Z => n1762);
   U1755 : AN2I port map( A => n1778, B => n1779, Z => n1773);
   U1762 : AN2I port map( A => n1778, B => n1781, Z => n1780);
   U1770 : AN2I port map( A => n1778, B => n1787, Z => n1786);
   U1777 : AN2I port map( A => n1778, B => n1789, Z => n1788);
   U1778 : NR2I port map( A => n8296, B => n8295, Z => n1778);
   U1786 : AN2I port map( A => n1797, B => n1779, Z => n1796);
   U1793 : AN2I port map( A => n1797, B => n1781, Z => n1798);
   U1801 : AN2I port map( A => n1797, B => n1787, Z => n1803);
   U1808 : AN2I port map( A => n1797, B => n1789, Z => n1804);
   U1809 : NR2I port map( A => n1805, B => n8296, Z => n1797);
   U1819 : AN2I port map( A => n1779, B => n1816, Z => n1815);
   U1826 : AN2I port map( A => n1781, B => n1816, Z => n1817);
   U1834 : AN2I port map( A => n1787, B => n1816, Z => n1822);
   U1841 : AN2I port map( A => n1789, B => n1816, Z => n1823);
   U1842 : NR2I port map( A => n1806, B => n8295, Z => n1816);
   U1851 : AN2I port map( A => n1829, B => n1779, Z => n1828);
   U1852 : NR2I port map( A => n8293, B => n8294, Z => n1779);
   U1859 : AN2I port map( A => n1829, B => n1781, Z => n1832);
   U1860 : NR2I port map( A => n1833, B => n8294, Z => n1781);
   U1869 : AN2I port map( A => n1829, B => n1787, Z => n1839);
   U1870 : NR2I port map( A => n1834, B => n8293, Z => n1787);
   U1874 : NR2I port map( A => n8292, B => n8291, Z => n1774);
   U1876 : NR2I port map( A => n1843, B => n8292, Z => n1775);
   U1880 : NR2I port map( A => n1844, B => n8291, Z => n1776);
   U1883 : NR2I port map( A => n1843, B => n1844, Z => n1777);
   U1886 : AN2I port map( A => n1829, B => n1789, Z => n1840);
   U1887 : NR2I port map( A => n1834, B => n1833, Z => n1789);
   U1890 : NR2I port map( A => n1805, B => n1806, Z => n1829);
   U1896 : AO1P port map( A => n8264, B => n1853, C => n1854, D => n1855, Z => 
                           n1851);
   U1899 : AO1P port map( A => n2005, B => n8237, C => n1866, D => n1867, Z => 
                           n1850);
   U1903 : AO1P port map( A => n2005, B => n1876, C => n1877, D => n1878, Z => 
                           n1875);
   U1905 : ND2I port map( A => n1881, B => n1857, Z => n1876);
   U1908 : ND2I port map( A => n381, B => n1890, Z => n1846);
   U1916 : ND2I port map( A => n276, B => n1915, Z => n1914);
   U1918 : NR2I port map( A => n8252, B => n8233, Z => n1917);
   U1926 : NR2I port map( A => n1936, B => n1937, Z => n1912);
   U1927 : NR2I port map( A => n2262, B => n1938, Z => n1878);
   U1932 : AO1P port map( A => n2085, B => n1948, C => n1949, D => n1950, Z => 
                           n1946);
   U1934 : ND2I port map( A => n8239, B => n8269, Z => n1952);
   U1936 : ND2I port map( A => n1957, B => n1958, Z => n1948);
   U1938 : NR2I port map( A => n8230, B => n8253, Z => n1884);
   U1940 : AO1P port map( A => n1963, B => n267, C => n1965, D => n1966, Z => 
                           n1962);
   U1941 : NR2I port map( A => n1967, B => n1968, Z => n1966);
   U1943 : AO1P port map( A => n1937, B => n267, C => n1970, D => n1971, Z => 
                           n1961);
   U1945 : ND2I port map( A => n1934, B => n1973, Z => n1972);
   U1951 : ND2I port map( A => n2183, B => n2234, Z => n1984);
   U1955 : ND2I port map( A => n1994, B => n1995, Z => n1991);
   U1957 : ND2I port map( A => n1996, B => n2214, Z => n1977);
   U1960 : ND2I port map( A => n1968, B => n1958, Z => n2003);
   U1961 : NR2I port map( A => n8251, B => n8247, Z => n2002);
   U1972 : NR2I port map( A => n376, B => n8230, Z => n1858);
   U1974 : AN2I port map( A => n2026, B => n2022, Z => n2025);
   U1975 : ND2I port map( A => n8226, B => n369, Z => n2022);
   U1991 : ND2I port map( A => n2189, B => n1969, Z => n2048);
   U1993 : ND2I port map( A => n1957, B => n1857, Z => n1853);
   U1998 : NR2I port map( A => n8231, B => n8223, Z => n1886);
   U2003 : NR2I port map( A => n8229, B => n2062, Z => n2061);
   U2007 : AO1P port map( A => n2072, B => n2073, C => n2074, D => n2075, Z => 
                           n2071);
   U2010 : ND2I port map( A => n2174, B => n2206, Z => n1900);
   U2026 : NR2I port map( A => n2102, B => n2103, Z => n2101);
   U2029 : NR2I port map( A => n2105, B => n2106, Z => n2100);
   U2034 : AO1P port map( A => n378, B => n2110, C => n8273, D => n2112, Z => 
                           n2097);
   U2037 : NR2I port map( A => n2115, B => n2183, Z => n2096);
   U2040 : AO1P port map( A => n8264, B => n2169, C => n2122, D => n2123, Z => 
                           n2121);
   U2042 : NR2I port map( A => n8264, B => n368, Z => n2124);
   U2046 : ND2I port map( A => n1994, B => n2127, Z => n1980);
   U2053 : NR2I port map( A => n8223, B => n8232, Z => n2135);
   U2054 : ND2I port map( A => n2138, B => n2139, Z => n2131);
   U2058 : AO1P port map( A => n2141, B => n2142, C => n2143, D => n2214, Z => 
                           n2129);
   U2061 : ND2I port map( A => n1963, B => n2085, Z => n2145);
   U2067 : NR2I port map( A => n8231, B => n2078, Z => n2149);
   U2068 : NR2I port map( A => n8224, B => n1879, Z => n2032);
   U2073 : ND2I port map( A => n2035, B => n2206, Z => n2056);
   U2077 : AO1P port map( A => n2005, B => n1993, C => n2159, D => n2160, Z => 
                           n2158);
   U2083 : ND2I port map( A => n1956, B => n2104, Z => n1993);
   U2085 : NR2I port map( A => n8229, B => n2078, Z => n2079);
   U2086 : NR2I port map( A => n8244, B => n2078, Z => n1870);
   U2088 : ND2I port map( A => n8274, B => n2214, Z => n2013);
   U2090 : ND2I port map( A => n2165, B => n8234, Z => n2164);
   U2096 : NR2I port map( A => n1937, B => n8255, Z => n2114);
   U2097 : NR2I port map( A => n2169, B => n1888, Z => n1937);
   U2100 : ND2I port map( A => n1958, B => n2127, Z => n2173);
   U2101 : ND2I port map( A => n8251, B => n2027, Z => n1958);
   U2104 : NR2I port map( A => n8235, B => n1880, Z => n2170);
   U2107 : AO1P port map( A => n2180, B => n2062, C => n2181, D => n2182, Z => 
                           n2179);
   U2110 : ND2I port map( A => n1934, B => n2287, Z => n2054);
   U2111 : EOI port map( A => n276, B => n2027, Z => n2062);
   U2112 : NR2I port map( A => n8229, B => n8267, Z => n2180);
   U2113 : AO1P port map( A => n8265, B => n8246, C => n2184, D => n1929, Z => 
                           n2178);
   U2114 : NR2I port map( A => n1881, B => n1967, Z => n1929);
   U2118 : ND2I port map( A => n1957, B => n2011, Z => n2186);
   U2119 : ND2I port map( A => n2115, B => n2187, Z => n1916);
   U2120 : AO1P port map( A => n8251, B => n2005, C => n8273, D => n2188, Z => 
                           n2175);
   U2129 : NR2I port map( A => n8235, B => n8231, Z => n2201);
   U2131 : ND2I port map( A => n2027, B => n1973, Z => n1857);
   U2133 : NR2I port map( A => n2035, B => n2206, Z => n2046);
   U2135 : NR2I port map( A => n8224, B => n8255, Z => n2008);
   U2138 : ND2I port map( A => n1925, B => n2214, Z => n1867);
   U2142 : ND2I port map( A => n8259, B => n267, Z => n2026);
   U2144 : ND2I port map( A => n2011, B => n2169, Z => n1934);
   U2145 : ND2I port map( A => n8229, B => n2169, Z => n2127);
   U2148 : NR2I port map( A => n8251, B => n2078, Z => n2137);
   U2150 : NR2I port map( A => n2214, B => n8273, Z => n1941);
   U2152 : NR2I port map( A => n8239, B => n8235, Z => n2053);
   U2154 : ND2I port map( A => n377, B => n2169, Z => n2104);
   U2155 : NR2I port map( A => n1879, B => n8259, Z => n2144);
   U2159 : ND2I port map( A => n1968, B => n2093, Z => n2031);
   U2162 : ND2I port map( A => n2027, B => n2136, Z => n1994);
   U2167 : ND2I port map( A => n1938, B => n2060, Z => n1928);
   U2169 : ND2I port map( A => n2218, B => n2214, Z => n2207);
   U2173 : ND2I port map( A => n8243, B => n2169, Z => n1995);
   U2174 : ND2I port map( A => n2082, B => n1938, Z => n2223);
   U2182 : NR2I port map( A => n8250, B => n8253, Z => n1860);
   U2186 : ND2I port map( A => v_SUB_WORD_7_port, B => n8165, Z => n2226);
   U2188 : NR2I port map( A => n2229, B => n2230, Z => n2228);
   U2190 : ND2I port map( A => n381, B => n274, Z => n1990);
   U2192 : ND2I port map( A => n1975, B => n8263, Z => n2232);
   U2193 : NR2I port map( A => n1936, B => n8245, Z => n1975);
   U2194 : ND2I port map( A => n1957, B => n2115, Z => n2210);
   U2196 : ND2I port map( A => n381, B => n2206, Z => n1983);
   U2202 : ND2I port map( A => n8142, B => n2237, Z => n1894);
   U2203 : AO1P port map( A => n2238, B => n2206, C => n2239, D => n2240, Z => 
                           n2227);
   U2205 : ND2I port map( A => n8246, B => n1922, Z => n2010);
   U2210 : EOI port map( A => n8267, B => n2169, Z => n2072);
   U2211 : NR2I port map( A => n2206, B => n8267, Z => n2040);
   U2213 : ND2I port map( A => n8251, B => n2169, Z => n2134);
   U2218 : ND2I port map( A => n2082, B => n1922, Z => n2244);
   U2219 : ND2I port map( A => n8229, B => n2027, Z => n1922);
   U2221 : ND2I port map( A => n8258, B => n267, Z => n2233);
   U2222 : NR2I port map( A => n8259, B => n8255, Z => n2242);
   U2225 : NR2I port map( A => n2237, B => n8166, Z => n1925);
   U2226 : ND2I port map( A => n2245, B => n2246, Z => n2237);
   U2231 : AO1P port map( A => n2128, B => n2253, C => n2254, D => n2255, Z => 
                           n2252);
   U2233 : ND2I port map( A => n8265, B => n274, Z => n1859);
   U2234 : ND2I port map( A => n2027, B => n2147, Z => n1938);
   U2236 : ND2I port map( A => n8262, B => n1957, Z => n2257);
   U2237 : ND2I port map( A => n370, B => n274, Z => n1871);
   U2240 : ND2I port map( A => n2027, B => n1888, Z => n1956);
   U2242 : ND2I port map( A => n8267, B => n2206, Z => n2162);
   U2243 : NR2I port map( A => n1936, B => n2028, Z => n1923);
   U2244 : NR2I port map( A => n1879, B => n1880, Z => n2128);
   U2245 : NR2I port map( A => n2147, B => n2027, Z => n1879);
   U2247 : NR2I port map( A => n8255, B => n8232, Z => n2109);
   U2249 : ND2I port map( A => n8233, B => n2027, Z => n2088);
   U2252 : ND2I port map( A => n2169, B => n2065, Z => n1968);
   U2253 : ND2I port map( A => n8263, B => n273, Z => n1861);
   U2254 : ND2I port map( A => n8246, B => n2115, Z => n2083);
   U2255 : ND2I port map( A => n2027, B => n2065, Z => n2115);
   U2257 : ND2I port map( A => n267, B => n274, Z => n1856);
   U2258 : NR2I port map( A => n8256, B => n2028, Z => n1872);
   U2261 : ND2I port map( A => n1957, B => n2147, Z => n2259);
   U2262 : ND2I port map( A => n267, B => n2206, Z => n1869);
   U2264 : NR2I port map( A => n8256, B => n1880, Z => n2107);
   U2265 : NR2I port map( A => n2011, B => n2169, Z => n1880);
   U2267 : ND2I port map( A => n8257, B => n2169, Z => n1881);
   U2270 : NR2I port map( A => n2028, B => n8258, Z => n1963);
   U2272 : ND2I port map( A => n2169, B => n1888, Z => n2060);
   U2274 : AO1P port map( A => n1868, B => n2005, C => n2214, D => n2260, Z => 
                           n2248);
   U2275 : AO1P port map( A => n267, B => n2065, C => n2261, D => n8225, Z => 
                           n2260);
   U2279 : ND2I port map( A => n8267, B => n2174, Z => n1969);
   U2280 : ND2I port map( A => n1882, B => n8246, Z => n2213);
   U2282 : NR2I port map( A => n2011, B => n2027, Z => n1936);
   U2283 : ND2I port map( A => n2027, B => n8243, Z => n1882);
   U2286 : ND2I port map( A => n2027, B => n2011, Z => n2093);
   U2296 : ND2I port map( A => n2169, B => n1973, Z => n2082);
   U2297 : ND2I port map( A => n8243, B => n1888, Z => n1973);
   U2299 : ND2I port map( A => n8267, B => n276, Z => n1924);
   U2301 : ND2I port map( A => n2264, B => n2265, Z => n1997);
   U2305 : ND2I port map( A => n370, B => n2206, Z => n1951);
   U2306 : ND2I port map( A => n2266, B => n2267, Z => n1911);
   U2310 : ND2I port map( A => n276, B => n2035, Z => n1935);
   U2315 : ND2I port map( A => n2270, B => n2271, Z => n1905);
   U2320 : ND2I port map( A => n2169, B => n2136, Z => n2187);
   U2322 : ND2I port map( A => n8243, B => n8257, Z => n2147);
   U2325 : ND2I port map( A => n2272, B => n2273, Z => n1927);
   U2329 : ND2I port map( A => n2065, B => n1888, Z => n2011);
   U2333 : ND2I port map( A => n2276, B => n2277, Z => n2065);
   U2336 : ND2I port map( A => v_CALCULATION_CNTR_1_port, B => n1985, Z => 
                           n2280);
   U2338 : ND2I port map( A => n8289, B => n367, Z => n2282);
   U2340 : ND2I port map( A => n2305, B => n2283, Z => n2278);
   U2343 : ND2I port map( A => n2285, B => n2286, Z => n2247);
   U2346 : NR2I port map( A => n231, B => n175, Z => n166);
   U2349 : ND2I port map( A => v_CALCULATION_CNTR_0_port, B => 
                           v_CALCULATION_CNTR_1_port, Z => n2281);
   U2353 : ND2I port map( A => VALID_KEY_I, B => n8143, Z => n336);
   U4469 : ND2I port map( A => n6638, B => n2467, Z => n2462);
   U4580 : ND2I port map( A => n8290, B => n8280, Z => n68);
   U4581 : NR2I port map( A => n2305, B => n367, Z => n2479);
   U4583 : ND2I port map( A => n2033, B => n8280, Z => n2285);
   U4585 : ND2I port map( A => n367, B => n1985, Z => n259);
   U4586 : NR2I port map( A => n236, B => n365, Z => n2284);
   U4595 : NR2I port map( A => n8297, B => n6638, Z => n2469);
   U4597 : NR2I port map( A => n8164, B => n2491, Z => n2467);
   U4627 : NR2I port map( A => n8143, B => RESET_I, Z => n2483);
   U4628 : NR2I port map( A => n269, B => n1903, Z => KEY_EXP_O(9));
   U4630 : NR2I port map( A => n269, B => n394, Z => KEY_EXP_O(8));
   U4632 : NR2I port map( A => n269, B => n354, Z => KEY_EXP_O(7));
   U4634 : NR2I port map( A => n269, B => n393, Z => KEY_EXP_O(6));
   U4636 : NR2I port map( A => n269, B => n382, Z => KEY_EXP_O(5));
   U4638 : NR2I port map( A => n269, B => n1630, Z => KEY_EXP_O(4));
   U4640 : NR2I port map( A => n2306, B => n1586, Z => KEY_EXP_O(3));
   U4642 : NR2I port map( A => n269, B => n1498, Z => KEY_EXP_O(31));
   U4644 : NR2I port map( A => n269, B => n353, Z => KEY_EXP_O(30));
   U4646 : NR2I port map( A => n269, B => n403, Z => KEY_EXP_O(2));
   U4648 : NR2I port map( A => n269, B => n392, Z => KEY_EXP_O(29));
   U4650 : NR2I port map( A => n2306, B => n1897, Z => KEY_EXP_O(28));
   U4652 : NR2I port map( A => n2306, B => n357, Z => KEY_EXP_O(27));
   U4654 : NR2I port map( A => n269, B => n391, Z => KEY_EXP_O(26));
   U4656 : NR2I port map( A => n2306, B => n1454, Z => KEY_EXP_O(25));
   U4658 : NR2I port map( A => n2306, B => n355, Z => KEY_EXP_O(24));
   U4660 : NR2I port map( A => n2306, B => n390, Z => KEY_EXP_O(23));
   U4662 : NR2I port map( A => n2306, B => n352, Z => KEY_EXP_O(22));
   U4664 : NR2I port map( A => n2306, B => n351, Z => KEY_EXP_O(21));
   U4666 : NR2I port map( A => n2306, B => n1906, Z => KEY_EXP_O(20));
   U4668 : NR2I port map( A => n2306, B => n1542, Z => KEY_EXP_O(1));
   U4670 : NR2I port map( A => n2306, B => n1367, Z => KEY_EXP_O(19));
   U4672 : NR2I port map( A => n2306, B => n389, Z => KEY_EXP_O(18));
   U4674 : NR2I port map( A => n2306, B => n1889, Z => KEY_EXP_O(17));
   U4676 : NR2I port map( A => n269, B => n388, Z => KEY_EXP_O(16));
   U4678 : NR2I port map( A => n2306, B => n387, Z => KEY_EXP_O(15));
   U4680 : NR2I port map( A => n269, B => n339, Z => KEY_EXP_O(14));
   U4682 : NR2I port map( A => n2306, B => n380, Z => KEY_EXP_O(13));
   U4684 : NR2I port map( A => n2306, B => n1904, Z => KEY_EXP_O(12));
   U4686 : NR2I port map( A => n2306, B => n356, Z => KEY_EXP_O(11));
   U4688 : NR2I port map( A => n2306, B => n327, Z => KEY_EXP_O(10));
   U4690 : NR2I port map( A => n269, B => n1887, Z => KEY_EXP_O(0));
   U3 : AO2 port map( A => v_TEMP_VECTOR_29_port, B => n2166, C => 
                           v_TEMP_VECTOR_21_port, D => n2168, Z => n2267);
   U4 : IVDAP port map( A => n1856, Y => n2085, Z => n2256);
   U5 : AO2 port map( A => n1928, B => n2005, C => n2031, D => n2085, Z => 
                           n2030);
   U6 : AO7 port map( A => n8251, B => n2169, C => n1881, Z => n2007);
   U8 : IVI port map( A => n1869, Z => n8260);
   U9 : IVI port map( A => n1969, Z => n8265);
   U10 : AO3 port map( A => n1912, B => n1900, C => n1913, D => n1914, Z => 
                           n1895);
   U11 : NR3 port map( A => n1900, B => n2076, C => n1899, Z => n2075);
   U13 : NR4 port map( A => n2131, B => n2132, C => n381, D => n2133, Z => 
                           n2130);
   U14 : AO4 port map( A => n2200, B => n1916, C => n274, D => n1917, Z => 
                           n1915);
   U15 : AO2 port map( A => n8228, B => n368, C => n8261, D => n2077, Z => 
                           n2138);
   U16 : EON1 port map( A => n376, B => n2257, C => n2064, D => n294, Z => 
                           n2254);
   U18 : EO1 port map( A => n8250, B => n2040, C => n2080, D => n377, Z => 
                           n2241);
   U19 : ND2I port map( A => n8257, B => n2065, Z => n2077);
   U20 : AO2 port map( A => n2020, B => n2200, C => n273, D => n2021, Z => 
                           n2019);
   U21 : AO4 port map( A => n6642, B => n237, C => n2095, D => n239, Z => n6699
                           );
   U23 : AO4 port map( A => n6648, B => n260, C => n2092, D => n262, Z => n6707
                           );
   U24 : EON1 port map( A => n367, B => n8301, C => N1748, D => n2482, Z => 
                           n6652);
   U25 : AO3 port map( A => n8140, B => n1954, C => n1846, D => n1847, Z => 
                           n4581);
   U26 : AO2 port map( A => n8272, B => n1849, C => n1850, D => n1851, Z => 
                           n1847);
   U28 : AO2 port map( A => n1941, B => n1942, C => n8271, D => n1944, Z => 
                           n1940);
   U29 : AO2 port map( A => n8272, B => n2069, C => n4545, D => n8145, Z => 
                           n2068);
   U30 : AO3 port map( A => n2116, B => n2117, C => n2118, D => n2119, Z => 
                           n4585);
   U31 : AO2 port map( A => n2175, B => n2176, C => n8274, D => n2177, Z => 
                           n2153);
   U33 : ND4 port map( A => n8274, B => n2207, C => n2208, D => n2209, Z => 
                           n2192);
   U34 : AN2I port map( A => n2452, B => n2453, Z => n1);
   U35 : AN2I port map( A => n2454, B => n2453, Z => n2);
   U36 : AN2I port map( A => n2455, B => n2453, Z => n3);
   U38 : AN2I port map( A => n2456, B => n2453, Z => n4);
   U39 : AN2I port map( A => n2457, B => n2453, Z => n5);
   U42 : AN2I port map( A => n2458, B => n2453, Z => n6);
   U43 : AN2I port map( A => n2459, B => n2453, Z => n7);
   U44 : AN2I port map( A => n2460, B => n2453, Z => n8);
   U46 : AN2I port map( A => n2464, B => n2452, Z => n9);
   U47 : AN2I port map( A => n2464, B => n2454, Z => n10);
   U50 : AN2I port map( A => n2464, B => n2455, Z => n11);
   U51 : AN2I port map( A => n2464, B => n2456, Z => n12);
   U53 : AN2I port map( A => n2464, B => n2457, Z => n14);
   U54 : AN2I port map( A => n2464, B => n2458, Z => n22);
   U55 : AN2I port map( A => n2464, B => n2459, Z => n23);
   U56 : AN2I port map( A => n2464, B => n2460, Z => n28);
   U58 : AN2I port map( A => n2465, B => n2452, Z => n33);
   U59 : AN2I port map( A => n2465, B => n2454, Z => n38);
   U60 : AN2I port map( A => n2465, B => n2455, Z => n43);
   U61 : AN2I port map( A => n2465, B => n2456, Z => n48);
   U63 : AN2I port map( A => n2465, B => n2457, Z => n53);
   U64 : AN2I port map( A => n2465, B => n2458, Z => n59);
   U65 : AN2I port map( A => n2465, B => n2459, Z => n63);
   U66 : AN2I port map( A => n2465, B => n2460, Z => n69);
   U68 : AN2I port map( A => n2466, B => n2452, Z => n71);
   U69 : AN2I port map( A => n2466, B => n2454, Z => n72);
   U70 : AN2I port map( A => n2466, B => n2455, Z => n81);
   U71 : AN2I port map( A => n2466, B => n2456, Z => n109);
   U73 : AN2I port map( A => n2466, B => n2457, Z => n122);
   U74 : AN2I port map( A => n2466, B => n2458, Z => n150);
   U75 : AN2I port map( A => n2466, B => n2459, Z => n163);
   U76 : AN2I port map( A => n2466, B => n2460, Z => n169);
   U78 : AN2I port map( A => n2468, B => n2457, Z => n170);
   U79 : AN2I port map( A => n2468, B => n2458, Z => n171);
   U80 : AN2I port map( A => n2468, B => n2459, Z => n181);
   U81 : AN2I port map( A => n2468, B => n2460, Z => n182);
   U83 : AN2I port map( A => n2470, B => n2457, Z => n188);
   U84 : AN2I port map( A => n2470, B => n2458, Z => n196);
   U85 : AN2I port map( A => n2470, B => n2459, Z => n198);
   U86 : AN2I port map( A => n2470, B => n2460, Z => n204);
   U88 : AN2I port map( A => n2471, B => n2457, Z => n206);
   U89 : AN2I port map( A => n2471, B => n2458, Z => n213);
   U92 : AN2I port map( A => n2471, B => n2459, Z => n221);
   U93 : AN2I port map( A => n2471, B => n2460, Z => n224);
   U94 : AN2I port map( A => n2472, B => n2457, Z => n233);
   U96 : AN2I port map( A => n2472, B => n2458, Z => n234);
   U97 : AN2I port map( A => n2472, B => n2459, Z => n235);
   U100 : AN2I port map( A => n2472, B => n2460, Z => n238);
   U101 : AN2I port map( A => n2468, B => n2452, Z => n240);
   U102 : AN2I port map( A => n2468, B => n2454, Z => n241);
   U103 : AN2I port map( A => n2468, B => n2455, Z => n242);
   U104 : AN2I port map( A => n2468, B => n2456, Z => n243);
   U106 : AN2I port map( A => n2470, B => n2452, Z => n244);
   U107 : AN2I port map( A => n2470, B => n2454, Z => n247);
   U108 : AN2I port map( A => n2470, B => n2455, Z => n248);
   U109 : AN2I port map( A => n2470, B => n2456, Z => n251);
   U111 : AN2I port map( A => n2471, B => n2452, Z => n252);
   U112 : AN2I port map( A => n2471, B => n2454, Z => n254);
   U113 : AN2I port map( A => n2471, B => n2455, Z => n255);
   U114 : AN2I port map( A => n2471, B => n2456, Z => n256);
   U116 : AN2I port map( A => n2472, B => n2452, Z => n261);
   U117 : AN2I port map( A => n2472, B => n2454, Z => n263);
   U118 : AN2I port map( A => n2472, B => n2455, Z => n264);
   U119 : AN2I port map( A => n2472, B => n2456, Z => n265);
   U121 : NR3P port map( A => n358, B => n4548, C => n288, Z => n266);
   U122 : NR2P port map( A => n266, B => n2475, Z => n271);
   U123 : IVDA port map( A => n1911, Y => n273, Z => n2200);
   U124 : AN2I port map( A => n2011, B => n2147, Z => n297);
   U126 : IVDAP port map( A => n166, Y => n364, Z => n2140);
   U127 : IVDA port map( A => v_CALCULATION_CNTR_2_port, Y => n366, Z => n2305)
                           ;
   U128 : IVDA port map( A => n297, Y => n376, Z => n377);
   U129 : IVDA port map( A => n1859, Y => n378, Z => n2288);
   U131 : AN2I port map( A => n1780, B => n2293, Z => n404);
   U132 : AN2I port map( A => n1780, B => n2295, Z => n405);
   U133 : AN2I port map( A => n1780, B => n2294, Z => n406);
   U134 : AN2I port map( A => n1773, B => n2293, Z => n407);
   U136 : AN2I port map( A => n1788, B => n2293, Z => n408);
   U137 : AN2I port map( A => n1788, B => n2295, Z => n409);
   U140 : AN2I port map( A => n1788, B => n2294, Z => n410);
   U141 : AN2I port map( A => n1786, B => n2293, Z => n415);
   U142 : AN2I port map( A => n1798, B => n2293, Z => n416);
   U144 : AN2I port map( A => n1798, B => n2295, Z => n417);
   U145 : AN2I port map( A => n1798, B => n2294, Z => n418);
   U148 : AN2I port map( A => n1796, B => n2293, Z => n419);
   U150 : AN2I port map( A => n1804, B => n2293, Z => n420);
   U151 : AN2I port map( A => n1804, B => n2295, Z => n421);
   U153 : AN2I port map( A => n1804, B => n2294, Z => n422);
   U155 : AN2I port map( A => n1803, B => n2293, Z => n427);
   U157 : AN2I port map( A => n2293, B => n1817, Z => n428);
   U158 : AN2I port map( A => n2295, B => n1817, Z => n429);
   U159 : AN2I port map( A => n2294, B => n1817, Z => n430);
   U160 : AN2I port map( A => n1815, B => n2293, Z => n431);
   U162 : AN2I port map( A => n1823, B => n2293, Z => n432);
   U164 : AN2I port map( A => n1823, B => n2295, Z => n433);
   U165 : AN2I port map( A => n1823, B => n2294, Z => n434);
   U166 : AN2I port map( A => n1822, B => n2293, Z => n439);
   U168 : AN2I port map( A => n1832, B => n2293, Z => n440);
   U170 : AN2I port map( A => n1832, B => n2295, Z => n441);
   U172 : AN2I port map( A => n1832, B => n2294, Z => n442);
   U173 : AN2I port map( A => n1828, B => n2293, Z => n443);
   U174 : AN2I port map( A => n1840, B => n2293, Z => n444);
   U176 : AN2I port map( A => n1840, B => n2295, Z => n445);
   U178 : AN2I port map( A => n1840, B => n2294, Z => n446);
   U180 : AN2I port map( A => n1839, B => n2293, Z => n447);
   U181 : AN2I port map( A => n1773, B => n2295, Z => n491);
   U182 : AN2I port map( A => n1773, B => n2294, Z => n535);
   U184 : AN2I port map( A => n1786, B => n2295, Z => n579);
   U186 : AN2I port map( A => n1786, B => n2294, Z => n623);
   U188 : AN2I port map( A => n1796, B => n2295, Z => n667);
   U189 : AN2I port map( A => n1796, B => n2294, Z => n754);
   U190 : AN2I port map( A => n1803, B => n2295, Z => n798);
   U192 : AN2I port map( A => n1803, B => n2294, Z => n842);
   U194 : AN2I port map( A => n1815, B => n2295, Z => n929);
   U196 : AN2I port map( A => n1815, B => n2294, Z => n973);
   U198 : AN2I port map( A => n1822, B => n2295, Z => n1017);
   U199 : AN2I port map( A => n1822, B => n2294, Z => n1104);
   U201 : AN2I port map( A => n1828, B => n2295, Z => n1148);
   U208 : AN2I port map( A => n1828, B => n2294, Z => n1192);
   U209 : AN2I port map( A => n1839, B => n2295, Z => n1279);
   U212 : AN2I port map( A => n1839, B => n2294, Z => n1323);
   U213 : AN2I port map( A => n1780, B => n2292, Z => n1674);
   U219 : AN2I port map( A => n1773, B => n2292, Z => n1718);
   U220 : AN2I port map( A => n1788, B => n2292, Z => n1790);
   U221 : AN2I port map( A => n1786, B => n2292, Z => n1791);
   U222 : AN2I port map( A => n1798, B => n2292, Z => n1830);
   U223 : AN2I port map( A => n1796, B => n2292, Z => n1831);
   U224 : AN2I port map( A => n1804, B => n2292, Z => n1841);
   U225 : AN2I port map( A => n1803, B => n2292, Z => n1842);
   U226 : AN2I port map( A => n2292, B => n1817, Z => n1845);
   U227 : AN2I port map( A => n1815, B => n2292, Z => n1848);
   U228 : AN2I port map( A => n1823, B => n2292, Z => n1852);
   U229 : AN2I port map( A => n1822, B => n2292, Z => n1862);
   U230 : AN2I port map( A => n1832, B => n2292, Z => n1864);
   U231 : AN2I port map( A => n1828, B => n2292, Z => n1865);
   U232 : AN2I port map( A => n1840, B => n2292, Z => n1883);
   U233 : AN2I port map( A => n1839, B => n2292, Z => n1885);
   U234 : ENI port map( A => i_INTERN_ADDR_RD0_5_port, B => n8170, Z => n1919);
   U236 : ENI port map( A => i_SRAM_ADDR_WR0_5_port, B => n8174, Z => n1920);
   U238 : EOI port map( A => n8169, B => i_INTERN_ADDR_RD0_4_port, Z => n1932);
   U239 : EOI port map( A => n8173, B => i_SRAM_ADDR_WR0_4_port, Z => n1943);
   U240 : ENI port map( A => n8168, B => i_INTERN_ADDR_RD0_3_port, Z => n1947);
   U242 : ENI port map( A => n8172, B => i_SRAM_ADDR_WR0_3_port, Z => n1953);
   U243 : EOI port map( A => n8167, B => i_INTERN_ADDR_RD0_2_port, Z => n1986);
   U245 : EOI port map( A => n8171, B => i_SRAM_ADDR_WR0_2_port, Z => n1989);
   U246 : B2I port map( A => n112, Z1 => n_3123, Z2 => n2166);
   U247 : AO3 port map( A => n8140, B => n1955, C => n1939, D => n1940, Z => 
                           n4582);
   U248 : EO1 port map( A => n2037, B => n8236, C => n2137, D => n1861, Z => 
                           n2029);
   U249 : ND4 port map( A => n8274, B => n1977, C => n2059, D => n1979, Z => 
                           n1939);
   U250 : AO2 port map( A => n2248, B => n2249, C => n2250, D => n2214, Z => 
                           n2224);
   U251 : ND3 port map( A => n2289, B => n317, C => v_CALCULATION_CNTR_3_port, 
                           Z => n236);
   U252 : AO2 port map( A => v_TEMP_VECTOR_31_port, B => n2166, C => 
                           v_TEMP_VECTOR_23_port, D => n2168, Z => n2271);
   U253 : AN2I port map( A => n369, B => n2206, Z => n2005);
   U254 : B2I port map( A => n1911, Z1 => n274, Z2 => n2206);
   U255 : AN3 port map( A => n2006, B => n2125, C => n2009, Z => n2289);
   U257 : AN2I port map( A => n1957, B => n2093, Z => n2049);
   U258 : B2I port map( A => n1871, Z1 => n294, Z2 => n2279);
   U259 : AO3 port map( A => n8241, B => n2234, C => n1987, D => n1988, Z => 
                           n2059);
   U260 : AO1 port map( A => n369, B => n2088, C => n273, D => n2148, Z => 
                           n2142);
   U261 : AN3P port map( A => n375, B => n317, C => n2043, Z => n2283);
   U262 : NR3 port map( A => n2050, B => n2051, C => n2052, Z => n2012);
   U264 : AO3 port map( A => n381, B => n2227, C => n8274, D => n2228, Z => 
                           n2225);
   U265 : AO2 port map( A => v_TEMP_VECTOR_15_port, B => n364, C => 
                           v_TEMP_VECTOR_7_port, D => n2247, Z => n2270);
   U267 : B3IP port map( A => n1905, Z1 => n276, Z2 => n2174);
   U269 : IVDAP port map( A => n1927, Y => n2027, Z => n2169);
   U271 : NR2I port map( A => n236, B => n366, Z => n2033);
   U272 : ND2I port map( A => n8263, B => n2206, Z => n1863);
   U274 : IVI port map( A => n8267, Z => n2035);
   U276 : IVI port map( A => n1896, Z => n8267);
   U277 : IVDA port map( A => n1859, Y => n2037, Z => n2290);
   U278 : AO4 port map( A => n1879, B => n2256, C => n1880, D => n1869, Z => 
                           n1877);
   U280 : AO2 port map( A => n8262, B => n2007, C => n2008, D => n8261, Z => 
                           n1999);
   U281 : AO4 port map( A => n2017, B => n2018, C => n2019, D => n1894, Z => 
                           n2016);
   U284 : ND2I port map( A => n2169, B => n2077, Z => n1957);
   U285 : AO1P port map( A => n8223, B => n2040, C => n2087, D => n381, Z => 
                           n2086);
   U287 : AO6 port map( A => n2187, B => n2287, C => n8267, Z => n2076);
   U288 : IVI port map( A => n1956, Z => n8259);
   U289 : AO3 port map( A => n8140, B => n1959, C => n2192, D => n2193, Z => 
                           n4587);
   U290 : AO3 port map( A => n2012, B => n2013, C => n2014, D => n2015, Z => 
                           n4583);
   U291 : AO3 port map( A => n2163, B => n2164, C => n2214, D => n1925, Z => 
                           n2154);
   U294 : NR3P port map( A => v_CALCULATION_CNTR_7_port, B => 
                           v_CALCULATION_CNTR_6_port, C => 
                           v_CALCULATION_CNTR_5_port, Z => n2043);
   U295 : ND2I port map( A => n370, B => n1991, Z => n2045);
   U296 : ND2I port map( A => n8263, B => n1993, Z => n2055);
   U297 : AN2I port map( A => n2045, B => n2055, Z => n1987);
   U299 : B2I port map( A => n153, Z1 => n_3124, Z2 => n2168);
   U301 : OR2P port map( A => n1879, B => n306, Z => n2110);
   U302 : OR2P port map( A => n8259, B => n8230, Z => n2064);
   U303 : AO1 port map( A => n8265, B => n1928, C => n2216, D => n2217, Z => 
                           n2215);
   U304 : AO1 port map( A => n2040, B => n2041, C => n2042, D => n8222, Z => 
                           n2039);
   U305 : AO1 port map( A => n2005, B => n8240, C => n2126, D => n1867, Z => 
                           n2120);
   U306 : EON1 port map( A => n1958, B => n2288, C => n294, D => n2081, Z => 
                           n2036);
   U307 : OR2P port map( A => n1937, B => n8258, Z => n2081);
   U308 : AO1 port map( A => n2107, B => n378, C => n2202, D => n1867, Z => 
                           n2196);
   U309 : IVDA port map( A => n1938, Y => n306, Z => n2287);
   U310 : IVDA port map( A => n1861, Y => n368, Z => n2262);
   U311 : AO4 port map( A => n2109, B => n2279, C => n1872, D => n2262, Z => 
                           n2108);
   U312 : IVI port map( A => n8053, Z => n8055);
   U313 : IVI port map( A => n8033, Z => n8035);
   U314 : IVI port map( A => n8013, Z => n8015);
   U315 : IVI port map( A => n7993, Z => n7995);
   U316 : IVI port map( A => n7973, Z => n7975);
   U317 : IVI port map( A => n7953, Z => n7955);
   U318 : IVI port map( A => n7933, Z => n7935);
   U319 : IVI port map( A => n7913, Z => n7915);
   U320 : IVI port map( A => n7893, Z => n7895);
   U321 : IVI port map( A => n7873, Z => n7875);
   U322 : IVI port map( A => n7853, Z => n7855);
   U323 : IVI port map( A => n7833, Z => n7835);
   U324 : IVI port map( A => n7813, Z => n7815);
   U325 : IVI port map( A => n7793, Z => n7795);
   U326 : IVI port map( A => n7773, Z => n7775);
   U327 : IVI port map( A => n7753, Z => n7755);
   U328 : IVI port map( A => n7733, Z => n7735);
   U329 : IVI port map( A => n7713, Z => n7715);
   U330 : IVI port map( A => n7693, Z => n7695);
   U331 : IVI port map( A => n7673, Z => n7675);
   U332 : IVI port map( A => n7653, Z => n7655);
   U333 : IVI port map( A => n7633, Z => n7635);
   U334 : IVI port map( A => n7613, Z => n7615);
   U335 : IVI port map( A => n7593, Z => n7595);
   U336 : IVI port map( A => n7573, Z => n7575);
   U337 : IVI port map( A => n7553, Z => n7555);
   U339 : IVI port map( A => n7533, Z => n7535);
   U340 : IVI port map( A => n7513, Z => n7515);
   U341 : IVI port map( A => n7493, Z => n7495);
   U342 : IVI port map( A => n7473, Z => n7475);
   U343 : IVI port map( A => n7453, Z => n7455);
   U344 : IVI port map( A => n7413, Z => n7415);
   U345 : IVI port map( A => n7393, Z => n7395);
   U346 : IVI port map( A => n7373, Z => n7375);
   U347 : IVI port map( A => n7353, Z => n7355);
   U348 : IVI port map( A => n7333, Z => n7335);
   U349 : IVI port map( A => n7313, Z => n7315);
   U350 : IVI port map( A => n7293, Z => n7295);
   U351 : IVI port map( A => n7253, Z => n7255);
   U352 : IVI port map( A => n7233, Z => n7235);
   U353 : IVI port map( A => n7213, Z => n7215);
   U354 : IVI port map( A => n7193, Z => n7195);
   U355 : IVI port map( A => n7173, Z => n7175);
   U357 : IVI port map( A => n7153, Z => n7155);
   U358 : IVI port map( A => n7133, Z => n7135);
   U359 : IVI port map( A => n7093, Z => n7095);
   U360 : IVI port map( A => n7073, Z => n7075);
   U361 : IVI port map( A => n7053, Z => n7055);
   U362 : IVI port map( A => n7033, Z => n7035);
   U363 : IVI port map( A => n7013, Z => n7015);
   U364 : IVI port map( A => n6993, Z => n6995);
   U365 : IVI port map( A => n6973, Z => n6975);
   U366 : IVI port map( A => n6933, Z => n6935);
   U367 : IVI port map( A => n6913, Z => n6915);
   U368 : IVI port map( A => n6893, Z => n6895);
   U369 : IVI port map( A => n6873, Z => n6875);
   U370 : IVI port map( A => n6853, Z => n6855);
   U371 : IVI port map( A => n6833, Z => n6835);
   U372 : IVI port map( A => n6813, Z => n6815);
   U373 : IVI port map( A => n8053, Z => n8054);
   U374 : IVI port map( A => n8033, Z => n8034);
   U375 : IVI port map( A => n8013, Z => n8014);
   U376 : IVI port map( A => n7993, Z => n7994);
   U378 : IVI port map( A => n7973, Z => n7974);
   U379 : IVI port map( A => n7953, Z => n7954);
   U380 : IVI port map( A => n7933, Z => n7934);
   U381 : IVI port map( A => n7913, Z => n7914);
   U383 : IVI port map( A => n7893, Z => n7894);
   U384 : IVI port map( A => n7873, Z => n7874);
   U385 : IVI port map( A => n7853, Z => n7854);
   U386 : IVI port map( A => n7833, Z => n7834);
   U387 : IVI port map( A => n7813, Z => n7814);
   U388 : IVI port map( A => n7793, Z => n7794);
   U389 : IVI port map( A => n7773, Z => n7774);
   U390 : IVI port map( A => n7753, Z => n7754);
   U391 : IVI port map( A => n7733, Z => n7734);
   U392 : IVI port map( A => n7713, Z => n7714);
   U393 : IVI port map( A => n7693, Z => n7694);
   U394 : IVI port map( A => n7673, Z => n7674);
   U395 : IVI port map( A => n7653, Z => n7654);
   U396 : IVI port map( A => n7633, Z => n7634);
   U397 : IVI port map( A => n7613, Z => n7614);
   U398 : IVI port map( A => n7593, Z => n7594);
   U399 : IVI port map( A => n7573, Z => n7574);
   U400 : IVI port map( A => n7553, Z => n7554);
   U401 : IVI port map( A => n7533, Z => n7534);
   U402 : IVI port map( A => n7513, Z => n7514);
   U403 : IVI port map( A => n7493, Z => n7494);
   U404 : IVI port map( A => n7473, Z => n7474);
   U405 : IVI port map( A => n7453, Z => n7454);
   U406 : IVI port map( A => n7413, Z => n7414);
   U407 : IVI port map( A => n7393, Z => n7394);
   U408 : IVI port map( A => n7373, Z => n7374);
   U409 : IVI port map( A => n7353, Z => n7354);
   U410 : IVI port map( A => n7333, Z => n7334);
   U411 : IVI port map( A => n7313, Z => n7314);
   U412 : IVI port map( A => n7293, Z => n7294);
   U413 : IVI port map( A => n7253, Z => n7254);
   U414 : IVI port map( A => n7233, Z => n7234);
   U415 : IVI port map( A => n7213, Z => n7214);
   U416 : IVI port map( A => n7193, Z => n7194);
   U417 : IVI port map( A => n7173, Z => n7174);
   U418 : IVI port map( A => n7153, Z => n7154);
   U419 : IVI port map( A => n7133, Z => n7134);
   U420 : IVI port map( A => n7093, Z => n7094);
   U421 : IVI port map( A => n7073, Z => n7074);
   U422 : IVI port map( A => n7053, Z => n7054);
   U423 : IVI port map( A => n7033, Z => n7034);
   U424 : IVI port map( A => n7013, Z => n7014);
   U425 : IVI port map( A => n6993, Z => n6994);
   U427 : IVI port map( A => n6973, Z => n6974);
   U428 : IVI port map( A => n6933, Z => n6934);
   U429 : IVI port map( A => n6913, Z => n6914);
   U430 : IVI port map( A => n6893, Z => n6894);
   U431 : IVI port map( A => n6873, Z => n6874);
   U432 : IVI port map( A => n6853, Z => n6854);
   U433 : IVI port map( A => n6833, Z => n6834);
   U434 : IVI port map( A => n6813, Z => n6814);
   U435 : IVI port map( A => n7433, Z => n7435);
   U436 : IVI port map( A => n7273, Z => n7275);
   U437 : IVI port map( A => n7113, Z => n7115);
   U438 : IVI port map( A => n6953, Z => n6955);
   U439 : IVI port map( A => n6793, Z => n6795);
   U440 : IVI port map( A => n7433, Z => n7434);
   U441 : IVI port map( A => n7273, Z => n7274);
   U442 : IVI port map( A => n7113, Z => n7114);
   U443 : IVI port map( A => n6953, Z => n6954);
   U444 : IVI port map( A => n6793, Z => n6794);
   U445 : IVI port map( A => n8165, Z => n8141);
   U446 : IVI port map( A => n8164, Z => n8140);
   U447 : IVI port map( A => n8165, Z => n8142);
   U448 : NR2I port map( A => n2027, B => n8233, Z => n2078);
   U449 : NR2I port map( A => n8244, B => n8236, Z => n1868);
   U450 : IVI port map( A => n1931, Z => n8264);
   U451 : IVI port map( A => n1863, Z => n8262);
   U452 : AO3 port map( A => n2144, B => n2290, C => n2145, D => n2146, Z => 
                           n2143);
   U453 : AO3 port map( A => n1872, B => n1951, C => n2251, D => n2252, Z => 
                           n2250);
   U454 : AO6 port map( A => n1881, B => n1938, C => n2290, Z => n2255);
   U455 : IVI port map( A => n2187, Z => n8236);
   U456 : EON1 port map( A => n1931, B => n8251, C => n1933, D => n1934, Z => 
                           n1930);
   U457 : AO7 port map( A => n1912, B => n2189, C => n2279, Z => n1933);
   U458 : IVI port map( A => n1957, Z => n8252);
   U459 : AO4 port map( A => n1860, B => n2262, C => n377, D => n1863, Z => 
                           n1854);
   U460 : AO3 port map( A => n2170, B => n1863, C => n2171, D => n2172, Z => 
                           n2163);
   U461 : AO6 port map( A => n1963, B => n8262, C => n2258, Z => n2249);
   U462 : AO2 port map( A => n8265, B => n2244, C => n8224, D => n369, Z => 
                           n2243);
   U463 : AO6 port map( A => n8242, B => n8265, C => n1990, Z => n1988);
   U464 : AO2 port map( A => n369, B => n2213, C => n8239, D => n8265, Z => 
                           n2211);
   U465 : IVDA port map( A => n1924, Y => n267, Z => n2234);
   U466 : IVDA port map( A => n80, Y => n_3125, Z => n2302);
   U467 : IVDA port map( A => n21, Y => n_3126, Z => n2304);
   U468 : IVDA port map( A => n80, Y => n_3127, Z => n2301);
   U469 : IVDA port map( A => n21, Y => n_3128, Z => n2303);
   U471 : AO6 port map( A => n8229, B => n8265, C => n1983, Z => n1982);
   U472 : AO6 port map( A => n267, B => n2031, C => n1983, Z => n2212);
   U473 : AN2I port map( A => n297, B => n2027, Z => n2028);
   U474 : ND2I port map( A => n8265, B => n2206, Z => n1931);
   U475 : AO4 port map( A => n1963, B => n8268, C => n2201, D => n1951, Z => 
                           n2199);
   U476 : AO4 port map( A => n2079, B => n2262, C => n8229, D => n2080, Z => 
                           n2074);
   U477 : NR3 port map( A => n273, B => n2096, C => n2113, Z => n2112);
   U478 : AO4 port map( A => n8251, B => n2234, C => n2049, D => n2191, Z => 
                           n2190);
   U479 : AO2 port map( A => n2005, B => n2144, C => n8262, D => n2053, Z => 
                           n2205);
   U480 : AO4 port map( A => n377, B => n2183, C => n1872, D => n1969, Z => 
                           n1965);
   U481 : EON1 port map( A => n2135, B => n1951, C => n2041, D => n8266, Z => 
                           n2132);
   U482 : AO4 port map( A => n1961, B => n2200, C => n273, D => n1962, Z => 
                           n1942);
   U483 : ND3 port map( A => n1925, B => n2029, C => n2030, Z => n2018);
   U484 : AO3 port map( A => n2287, B => n2056, C => n2057, D => n2058, Z => 
                           n2050);
   U485 : AO2 port map( A => n2046, B => n8250, C => n2005, D => n2060, Z => 
                           n2058);
   U486 : AO2 port map( A => n2061, B => n2040, C => n2062, D => n2063, Z => 
                           n2057);
   U487 : AO4 port map( A => n2178, B => n2206, C => n274, D => n2179, Z => 
                           n2177);
   U488 : AO3 port map( A => n8229, B => n2290, C => n2157, D => n2158, Z => 
                           n2156);
   U489 : IVI port map( A => n1967, Z => n8263);
   U490 : AO4 port map( A => n377, B => n2279, C => n2109, D => n1863, Z => 
                           n2122);
   U491 : AO2 port map( A => n8256, B => n2037, C => n8251, D => n8262, Z => 
                           n2139);
   U492 : AO7 port map( A => n2011, B => n2080, C => n2026, Z => n2204);
   U493 : AO7 port map( A => n8226, B => n1937, C => n8266, Z => n2161);
   U494 : AO2 port map( A => n8262, B => n2169, C => n2037, D => n1928, Z => 
                           n1926);
   U495 : AO7 port map( A => n2183, B => n2007, C => n2236, Z => n2235);
   U496 : AO7 port map( A => n232, B => n8162, C => n8286, Z => n172);
   U497 : IVDA port map( A => n1935, Y => n369, Z => n2183);
   U498 : AO4 port map( A => n2279, B => n1937, C => n2290, D => n1923, Z => 
                           n2089);
   U499 : AO7 port map( A => n66, B => n2166, C => n67, Z => n108);
   U500 : AO7 port map( A => n66, B => n62, C => n67, Z => n57);
   U501 : IVDA port map( A => n121, Y => n_3129, Z => n2300);
   U502 : OR3 port map( A => n2166, B => n8281, C => n8278, Z => n80);
   U503 : OR3 port map( A => n62, B => n8281, C => n8221, Z => n21);
   U504 : IVDA port map( A => n121, Y => n_3130, Z => n2299);
   U505 : IVI port map( A => n6732, Z => n6730);
   U506 : IVI port map( A => n6732, Z => n6729);
   U507 : IVI port map( A => n6732, Z => n6728);
   U508 : IVI port map( A => n6732, Z => n6727);
   U509 : IVI port map( A => n2402, Z => n2400);
   U510 : IVI port map( A => n2402, Z => n2399);
   U511 : IVI port map( A => n2402, Z => n2398);
   U512 : IVI port map( A => n2402, Z => n2397);
   U513 : IVI port map( A => n2354, Z => n2352);
   U515 : IVI port map( A => n2354, Z => n2351);
   U516 : IVI port map( A => n2354, Z => n2350);
   U517 : IVI port map( A => n2354, Z => n2349);
   U518 : IVI port map( A => n8062, Z => n8060);
   U519 : IVI port map( A => n8062, Z => n8059);
   U520 : IVI port map( A => n8062, Z => n8058);
   U521 : IVI port map( A => n8062, Z => n8057);
   U522 : IVI port map( A => n6726, Z => n6724);
   U523 : IVI port map( A => n6726, Z => n6723);
   U524 : IVI port map( A => n6726, Z => n6722);
   U525 : IVI port map( A => n6726, Z => n6721);
   U526 : IVI port map( A => n2396, Z => n2394);
   U527 : IVI port map( A => n2396, Z => n2393);
   U528 : IVI port map( A => n2396, Z => n2392);
   U529 : IVI port map( A => n2396, Z => n2391);
   U530 : IVI port map( A => n2348, Z => n2346);
   U531 : IVI port map( A => n2348, Z => n2345);
   U532 : IVI port map( A => n2348, Z => n2344);
   U533 : IVI port map( A => n2348, Z => n2343);
   U534 : IVI port map( A => n6776, Z => n6774);
   U535 : IVI port map( A => n6776, Z => n6773);
   U536 : IVI port map( A => n6776, Z => n6772);
   U537 : IVI port map( A => n6776, Z => n6771);
   U538 : IVI port map( A => n6720, Z => n6718);
   U539 : IVI port map( A => n6720, Z => n6717);
   U540 : IVI port map( A => n6720, Z => n6716);
   U541 : IVI port map( A => n6720, Z => n6658);
   U542 : IVI port map( A => n2390, Z => n2388);
   U543 : IVI port map( A => n2390, Z => n2387);
   U544 : IVI port map( A => n2390, Z => n2386);
   U545 : IVI port map( A => n2390, Z => n2385);
   U546 : IVI port map( A => n2342, Z => n2340);
   U547 : IVI port map( A => n2342, Z => n2339);
   U548 : IVI port map( A => n2342, Z => n2338);
   U549 : IVI port map( A => n2342, Z => n2337);
   U550 : IVI port map( A => n6770, Z => n6768);
   U551 : IVI port map( A => n6770, Z => n6767);
   U552 : IVI port map( A => n6770, Z => n6766);
   U553 : IVI port map( A => n6770, Z => n6765);
   U554 : IVI port map( A => n6657, Z => n6650);
   U555 : IVI port map( A => n6657, Z => n4543);
   U556 : IVI port map( A => n6657, Z => n4542);
   U557 : IVI port map( A => n6657, Z => n2490);
   U559 : IVI port map( A => n2384, Z => n2382);
   U560 : IVI port map( A => n2384, Z => n2381);
   U561 : IVI port map( A => n2384, Z => n2380);
   U562 : IVI port map( A => n2384, Z => n2379);
   U563 : IVI port map( A => n2336, Z => n2334);
   U564 : IVI port map( A => n2336, Z => n2333);
   U565 : IVI port map( A => n2336, Z => n2332);
   U566 : IVI port map( A => n2336, Z => n2331);
   U567 : IVI port map( A => n6764, Z => n6762);
   U568 : IVI port map( A => n6764, Z => n6761);
   U569 : IVI port map( A => n6764, Z => n6760);
   U570 : IVI port map( A => n6764, Z => n6759);
   U571 : IVI port map( A => n2481, Z => n2474);
   U572 : IVI port map( A => n2481, Z => n2473);
   U573 : IVI port map( A => n2481, Z => n2463);
   U574 : IVI port map( A => n2481, Z => n2461);
   U575 : IVI port map( A => n2378, Z => n2376);
   U576 : IVI port map( A => n2378, Z => n2375);
   U577 : IVI port map( A => n2378, Z => n2374);
   U578 : IVI port map( A => n2378, Z => n2373);
   U579 : IVI port map( A => n2330, Z => n2328);
   U580 : IVI port map( A => n2330, Z => n2327);
   U581 : IVI port map( A => n2330, Z => n2326);
   U582 : IVI port map( A => n2330, Z => n2325);
   U583 : IVI port map( A => n6758, Z => n6756);
   U584 : IVI port map( A => n6758, Z => n6755);
   U585 : IVI port map( A => n6758, Z => n6754);
   U586 : IVI port map( A => n6758, Z => n6753);
   U587 : IVI port map( A => n2420, Z => n2418);
   U588 : IVI port map( A => n2420, Z => n2417);
   U589 : IVI port map( A => n2420, Z => n2416);
   U590 : IVI port map( A => n2420, Z => n2415);
   U591 : IVI port map( A => n2372, Z => n2370);
   U592 : IVI port map( A => n2372, Z => n2369);
   U593 : IVI port map( A => n2372, Z => n2368);
   U594 : IVI port map( A => n2372, Z => n2367);
   U595 : IVI port map( A => n2324, Z => n2322);
   U596 : IVI port map( A => n2324, Z => n2321);
   U597 : IVI port map( A => n2324, Z => n2320);
   U598 : IVI port map( A => n2324, Z => n2319);
   U599 : IVI port map( A => n6752, Z => n6750);
   U600 : IVI port map( A => n6752, Z => n6747);
   U601 : IVI port map( A => n6752, Z => n6746);
   U603 : IVI port map( A => n6752, Z => n6745);
   U604 : IVI port map( A => n2414, Z => n2412);
   U605 : IVI port map( A => n2414, Z => n2411);
   U606 : IVI port map( A => n2414, Z => n2410);
   U607 : IVI port map( A => n2414, Z => n2409);
   U608 : IVI port map( A => n2366, Z => n2364);
   U609 : IVI port map( A => n2366, Z => n2363);
   U610 : IVI port map( A => n2366, Z => n2362);
   U611 : IVI port map( A => n2366, Z => n2361);
   U612 : IVI port map( A => n2318, Z => n2316);
   U613 : IVI port map( A => n2318, Z => n2315);
   U614 : IVI port map( A => n2318, Z => n2314);
   U615 : IVI port map( A => n2318, Z => n2313);
   U616 : IVI port map( A => n6744, Z => n6742);
   U617 : IVI port map( A => n6744, Z => n6741);
   U618 : IVI port map( A => n6744, Z => n6740);
   U619 : IVI port map( A => n6744, Z => n6739);
   U620 : IVI port map( A => n2408, Z => n2406);
   U621 : IVI port map( A => n2408, Z => n2405);
   U622 : IVI port map( A => n2408, Z => n2404);
   U623 : IVI port map( A => n2408, Z => n2403);
   U624 : IVI port map( A => n2360, Z => n2358);
   U625 : IVI port map( A => n2360, Z => n2357);
   U626 : IVI port map( A => n2360, Z => n2356);
   U627 : IVI port map( A => n2360, Z => n2355);
   U628 : IVI port map( A => n2312, Z => n2310);
   U629 : IVI port map( A => n2312, Z => n2309);
   U630 : IVI port map( A => n2312, Z => n2308);
   U631 : IVI port map( A => n2312, Z => n2307);
   U632 : IVI port map( A => n6738, Z => n6736);
   U633 : IVI port map( A => n6738, Z => n6735);
   U634 : IVI port map( A => n6738, Z => n6734);
   U635 : IVI port map( A => n6738, Z => n6733);
   U636 : IVDA port map( A => n1774, Y => n_3131, Z => n2295);
   U637 : ND2I port map( A => n1896, B => n2174, Z => n1967);
   U638 : AO2 port map( A => n8263, B => n2083, C => n2149, D => n8265, Z => 
                           n2141);
   U639 : AO4 port map( A => n276, B => n2137, C => n2114, D => n2174, Z => 
                           n2041);
   U640 : AO4 port map( A => n2281, B => n8288, C => n1985, D => n2282, Z => 
                           n112);
   U641 : AO7 port map( A => n8230, B => n2189, C => n274, Z => n2261);
   U642 : AO6 port map( A => n2028, B => n2035, C => n369, Z => n2191);
   U643 : AO4 port map( A => n1891, B => n1892, C => n1893, D => n1894, Z => 
                           n1890);
   U644 : AO3 port map( A => n1923, B => n2234, C => n1925, D => n1926, Z => 
                           n1892);
   U645 : AO2 port map( A => n2194, B => n2195, C => n2196, D => n2197, Z => 
                           n2193);
   U647 : ND3 port map( A => n1873, B => n1874, C => n1875, Z => n1849);
   U648 : AO2 port map( A => n8264, B => n1882, C => n8262, D => n1884, Z => 
                           n1874);
   U649 : ND4 port map( A => n1998, B => n1999, C => n2000, D => n2001, Z => 
                           n1996);
   U650 : AO2 port map( A => n8259, B => n368, C => n8228, D => n8264, Z => 
                           n2000);
   U651 : ND4 port map( A => n2219, B => n2220, C => n2221, D => n2222, Z => 
                           n2218);
   U652 : AO2 port map( A => n8264, B => n2223, C => n8223, D => n370, Z => 
                           n2222);
   U653 : AO4 port map( A => n2100, B => n2200, C => n273, D => n2101, Z => 
                           n2099);
   U654 : EO1 port map( A => n2047, B => n2048, C => n2048, D => n1870, Z => 
                           n2038);
   U655 : AO3 port map( A => n1899, B => n1900, C => n1901, D => n1902, Z => 
                           n1898);
   U656 : AO7 port map( A => n2090, B => n2091, C => n2200, Z => n2084);
   U657 : AO4 port map( A => n366, B => n68, C => n257, D => n258, Z => n157);
   U658 : AO7 port map( A => n66, B => n2168, C => n67, Z => n149);
   U659 : OR3 port map( A => n2168, B => n8281, C => n8276, Z => n121);
   U660 : EO1 port map( A => n2479, B => n8290, C => n68, D => n366, Z => n2478
                           );
   U661 : IVDA port map( A => n164, Y => n_3132, Z => n2297);
   U662 : AO4 port map( A => n2305, B => n68, C => n367, D => n70, Z => n62);
   U663 : AO7 port map( A => n268, B => n8163, C => n246, Z => n260);
   U664 : AO6 port map( A => n270, B => n366, C => n8281, Z => n268);
   U665 : IVDA port map( A => n1775, Y => n_3133, Z => n2294);
   U666 : IVDA port map( A => n1776, Y => n_3134, Z => n2293);
   U667 : IVDA port map( A => n1777, Y => n_3135, Z => n2292);
   U668 : AO4 port map( A => n8142, B => n394, C => n340, D => n8162, Z => 
                           n4549);
   U669 : ND4 port map( A => n395, B => n396, C => n397, D => n398, Z => n341);
   U670 : ND4 port map( A => n343, B => n344, C => n345, D => n346, Z => n342);
   U671 : AO4 port map( A => n8142, B => n388, C => n448, D => n8160, Z => 
                           n4550);
   U672 : ND4 port map( A => n471, B => n472, C => n473, D => n474, Z => n449);
   U673 : ND4 port map( A => n451, B => n452, C => n453, D => n454, Z => n450);
   U674 : AO4 port map( A => n8142, B => n355, C => n492, D => n8161, Z => 
                           n4551);
   U675 : ND4 port map( A => n515, B => n516, C => n517, D => n518, Z => n493);
   U676 : ND4 port map( A => n495, B => n496, C => n497, D => n498, Z => n494);
   U677 : AO4 port map( A => n8142, B => n1887, C => n536, D => n8159, Z => 
                           n4552);
   U678 : ND4 port map( A => n559, B => n560, C => n561, D => n562, Z => n537);
   U679 : ND4 port map( A => n539, B => n540, C => n541, D => n542, Z => n538);
   U680 : AO4 port map( A => n8142, B => n1903, C => n580, D => n8160, Z => 
                           n4553);
   U681 : ND4 port map( A => n603, B => n604, C => n605, D => n606, Z => n581);
   U682 : ND4 port map( A => n583, B => n584, C => n585, D => n586, Z => n582);
   U683 : AO4 port map( A => n8142, B => n1889, C => n624, D => n8158, Z => 
                           n4554);
   U684 : ND4 port map( A => n647, B => n648, C => n649, D => n650, Z => n625);
   U685 : ND4 port map( A => n627, B => n628, C => n629, D => n630, Z => n626);
   U686 : AO4 port map( A => n8142, B => n1454, C => n668, D => n8159, Z => 
                           n4555);
   U687 : ND4 port map( A => n691, B => n692, C => n693, D => n694, Z => n669);
   U688 : ND4 port map( A => n671, B => n672, C => n673, D => n674, Z => n670);
   U689 : AO4 port map( A => n8142, B => n1542, C => n711, D => n8157, Z => 
                           n4556);
   U691 : ND4 port map( A => n734, B => n735, C => n736, D => n737, Z => n712);
   U692 : ND4 port map( A => n714, B => n715, C => n716, D => n717, Z => n713);
   U693 : AO4 port map( A => n8142, B => n327, C => n755, D => n8158, Z => 
                           n4557);
   U694 : ND4 port map( A => n778, B => n779, C => n780, D => n781, Z => n756);
   U695 : ND4 port map( A => n758, B => n759, C => n760, D => n761, Z => n757);
   U696 : AO4 port map( A => n8141, B => n389, C => n799, D => n8156, Z => 
                           n4558);
   U697 : ND4 port map( A => n822, B => n823, C => n824, D => n825, Z => n800);
   U698 : ND4 port map( A => n802, B => n803, C => n804, D => n805, Z => n801);
   U699 : AO4 port map( A => n8141, B => n391, C => n843, D => n8157, Z => 
                           n4559);
   U700 : ND4 port map( A => n866, B => n867, C => n868, D => n869, Z => n844);
   U701 : ND4 port map( A => n846, B => n847, C => n848, D => n849, Z => n845);
   U702 : AO4 port map( A => n8141, B => n403, C => n886, D => n8155, Z => 
                           n4560);
   U703 : ND4 port map( A => n909, B => n910, C => n911, D => n912, Z => n887);
   U704 : ND4 port map( A => n889, B => n890, C => n891, D => n892, Z => n888);
   U705 : AO4 port map( A => n8141, B => n356, C => n930, D => n8156, Z => 
                           n4561);
   U706 : ND4 port map( A => n953, B => n954, C => n955, D => n956, Z => n931);
   U707 : ND4 port map( A => n933, B => n934, C => n935, D => n936, Z => n932);
   U708 : AO4 port map( A => n8141, B => n1367, C => n974, D => n8154, Z => 
                           n4562);
   U709 : ND4 port map( A => n997, B => n998, C => n999, D => n1000, Z => n975)
                           ;
   U710 : ND4 port map( A => n977, B => n978, C => n979, D => n980, Z => n976);
   U711 : AO4 port map( A => n8141, B => n357, C => n1018, D => n8155, Z => 
                           n4563);
   U712 : ND4 port map( A => n1041, B => n1042, C => n1043, D => n1044, Z => 
                           n1019);
   U713 : ND4 port map( A => n1021, B => n1022, C => n1023, D => n1024, Z => 
                           n1020);
   U714 : AO4 port map( A => n8141, B => n1586, C => n1061, D => n8154, Z => 
                           n4564);
   U715 : ND4 port map( A => n1084, B => n1085, C => n1086, D => n1087, Z => 
                           n1062);
   U716 : ND4 port map( A => n1064, B => n1065, C => n1066, D => n1067, Z => 
                           n1063);
   U717 : AO4 port map( A => n8141, B => n1904, C => n1105, D => n8153, Z => 
                           n4565);
   U718 : ND4 port map( A => n1128, B => n1129, C => n1130, D => n1131, Z => 
                           n1106);
   U719 : ND4 port map( A => n1108, B => n1109, C => n1110, D => n1111, Z => 
                           n1107);
   U720 : AO4 port map( A => n8141, B => n1906, C => n1149, D => n8153, Z => 
                           n4566);
   U721 : ND4 port map( A => n1172, B => n1173, C => n1174, D => n1175, Z => 
                           n1150);
   U722 : ND4 port map( A => n1152, B => n1153, C => n1154, D => n1155, Z => 
                           n1151);
   U723 : AO4 port map( A => n8141, B => n1897, C => n1193, D => n8152, Z => 
                           n4567);
   U724 : ND4 port map( A => n1216, B => n1217, C => n1218, D => n1219, Z => 
                           n1194);
   U725 : ND4 port map( A => n1196, B => n1197, C => n1198, D => n1199, Z => 
                           n1195);
   U726 : AO4 port map( A => n8141, B => n1630, C => n1236, D => n8152, Z => 
                           n4568);
   U727 : ND4 port map( A => n1259, B => n1260, C => n1261, D => n1262, Z => 
                           n1237);
   U728 : ND4 port map( A => n1239, B => n1240, C => n1241, D => n1242, Z => 
                           n1238);
   U729 : AO4 port map( A => n8141, B => n380, C => n1280, D => n8151, Z => 
                           n4569);
   U730 : ND4 port map( A => n1303, B => n1304, C => n1305, D => n1306, Z => 
                           n1281);
   U731 : ND4 port map( A => n1283, B => n1284, C => n1285, D => n1286, Z => 
                           n1282);
   U732 : AO4 port map( A => n8141, B => n351, C => n1324, D => n8151, Z => 
                           n4570);
   U733 : ND4 port map( A => n1347, B => n1348, C => n1349, D => n1350, Z => 
                           n1325);
   U735 : ND4 port map( A => n1327, B => n1328, C => n1329, D => n1330, Z => 
                           n1326);
   U736 : AO4 port map( A => n8140, B => n392, C => n1368, D => n8150, Z => 
                           n4571);
   U737 : ND4 port map( A => n1391, B => n1392, C => n1393, D => n1394, Z => 
                           n1369);
   U738 : ND4 port map( A => n1371, B => n1372, C => n1373, D => n1374, Z => 
                           n1370);
   U739 : AO4 port map( A => n8140, B => n382, C => n1411, D => n8150, Z => 
                           n4572);
   U740 : ND4 port map( A => n1434, B => n1435, C => n1436, D => n1437, Z => 
                           n1412);
   U741 : ND4 port map( A => n1414, B => n1415, C => n1416, D => n1417, Z => 
                           n1413);
   U742 : AO4 port map( A => n8140, B => n339, C => n1455, D => n8149, Z => 
                           n4573);
   U743 : ND4 port map( A => n1478, B => n1479, C => n1480, D => n1481, Z => 
                           n1456);
   U744 : ND4 port map( A => n1458, B => n1459, C => n1460, D => n1461, Z => 
                           n1457);
   U745 : AO4 port map( A => n8140, B => n352, C => n1499, D => n8149, Z => 
                           n4574);
   U746 : ND4 port map( A => n1522, B => n1523, C => n1524, D => n1525, Z => 
                           n1500);
   U747 : ND4 port map( A => n1502, B => n1503, C => n1504, D => n1505, Z => 
                           n1501);
   U748 : AO4 port map( A => n8140, B => n353, C => n1543, D => n8148, Z => 
                           n4575);
   U749 : ND4 port map( A => n1566, B => n1567, C => n1568, D => n1569, Z => 
                           n1544);
   U750 : ND4 port map( A => n1546, B => n1547, C => n1548, D => n1549, Z => 
                           n1545);
   U751 : AO4 port map( A => n8140, B => n393, C => n1587, D => n8148, Z => 
                           n4576);
   U752 : ND4 port map( A => n1610, B => n1611, C => n1612, D => n1613, Z => 
                           n1588);
   U753 : ND4 port map( A => n1590, B => n1591, C => n1592, D => n1593, Z => 
                           n1589);
   U754 : AO4 port map( A => n8141, B => n387, C => n1631, D => n8147, Z => 
                           n4577);
   U755 : ND4 port map( A => n1654, B => n1655, C => n1656, D => n1657, Z => 
                           n1632);
   U756 : ND4 port map( A => n1634, B => n1635, C => n1636, D => n1637, Z => 
                           n1633);
   U757 : AO4 port map( A => n8140, B => n390, C => n1675, D => n8147, Z => 
                           n4578);
   U758 : ND4 port map( A => n1698, B => n1699, C => n1700, D => n1701, Z => 
                           n1676);
   U759 : ND4 port map( A => n1678, B => n1679, C => n1680, D => n1681, Z => 
                           n1677);
   U760 : AO4 port map( A => n8140, B => n1498, C => n1719, D => n8146, Z => 
                           n4579);
   U761 : ND4 port map( A => n1742, B => n1743, C => n1744, D => n1745, Z => 
                           n1720);
   U762 : ND4 port map( A => n1722, B => n1723, C => n1724, D => n1725, Z => 
                           n1721);
   U763 : AO4 port map( A => n8140, B => n354, C => n1762, D => n8146, Z => 
                           n4580);
   U764 : ND4 port map( A => n1807, B => n1808, C => n1809, D => n1810, Z => 
                           n1763);
   U765 : ND4 port map( A => n1765, B => n1766, C => n1767, D => n1768, Z => 
                           n1764);
   U766 : NR4 port map( A => n1907, B => n65, C => n8285, D => n2483, Z => 
                           n2482);
   U767 : NR3 port map( A => i_SRAM_ADDR_WR0_3_port, B => n2462, C => 
                           i_SRAM_ADDR_WR0_4_port, Z => n2453);
   U768 : AO7 port map( A => n65, B => n290, C => n8283, Z => n287);
   U769 : AO7 port map( A => n8285, B => n155, C => n67, Z => n293);
   U770 : AO7 port map( A => n65, B => n190, C => n285, Z => n6712);
   U771 : AO2 port map( A => n207, B => n286, C => n287, D => n1918, Z => n285)
                           ;
   U772 : ND3 port map( A => n358, B => n288, C => n315, Z => n328);
   U773 : AO4 port map( A => n272, B => n1907, C => n8215, D => n275, Z => 
                           n6709);
   U774 : IVDA port map( A => n296, Y => n1909, Z => n2298);
   U775 : IVDA port map( A => n307, Y => n1910, Z => n2296);
   U776 : AO2 port map( A => v_TEMP_VECTOR_26_port, B => n2166, C => 
                           v_TEMP_VECTOR_18_port, D => n2168, Z => n2269);
   U777 : AO2 port map( A => v_TEMP_VECTOR_10_port, B => n364, C => 
                           v_TEMP_VECTOR_2_port, D => n2247, Z => n2268);
   U779 : AO2 port map( A => v_TEMP_VECTOR_27_port, B => n2166, C => 
                           v_TEMP_VECTOR_19_port, D => n2168, Z => n2275);
   U780 : AO2 port map( A => v_TEMP_VECTOR_11_port, B => n364, C => 
                           v_TEMP_VECTOR_3_port, D => n2247, Z => n2274);
   U781 : AO2 port map( A => v_TEMP_VECTOR_28_port, B => n2166, C => 
                           v_TEMP_VECTOR_20_port, D => n2168, Z => n2277);
   U782 : AO2 port map( A => v_TEMP_VECTOR_12_port, B => n364, C => 
                           v_TEMP_VECTOR_4_port, D => n2247, Z => n2276);
   U783 : AO4 port map( A => n2278, B => n259, C => n8288, D => n2280, Z => 
                           n153);
   U784 : AO2 port map( A => v_TEMP_VECTOR_25_port, B => n2166, C => 
                           v_TEMP_VECTOR_17_port, D => n2168, Z => n2273);
   U785 : AO3 port map( A => n274, B => n2038, C => n8271, D => n2039, Z => 
                           n2014);
   U786 : AO2 port map( A => n381, B => n2016, C => n4544, D => n8145, Z => 
                           n2015);
   U787 : AO3 port map( A => n2066, B => n2214, C => n2067, D => n2068, Z => 
                           n4584);
   U788 : ND4 port map( A => n1925, B => n2084, C => n8238, D => n2086, Z => 
                           n2067);
   U789 : AO2 port map( A => n2097, B => n2098, C => n8274, D => n2099, Z => 
                           n2066);
   U790 : AO3 port map( A => n2153, B => n2214, C => n2154, D => n2155, Z => 
                           n4586);
   U791 : AO2 port map( A => n8272, B => n2156, C => n4547, D => n8144, Z => 
                           n2155);
   U792 : AO3 port map( A => n2224, B => n8273, C => n2225, D => n2226, Z => 
                           n4588);
   U793 : AN3 port map( A => n367, B => v_CALCULATION_CNTR_0_port, C => n2284, 
                           Z => n231);
   U794 : ND4 port map( A => v_CALCULATION_CNTR_1_port, B => n2283, C => n1985,
                           D => n366, Z => n2286);
   U795 : AO7 port map( A => n1992, B => n172, C => n225, Z => n6695);
   U796 : AO2 port map( A => n2297, B => n226, C => v_KEY32_IN_0_port, D => 
                           n162, Z => n225);
   U797 : AO3 port map( A => n159, B => n216, C => n217, D => n218, Z => n6694)
                           ;
   U798 : AO2 port map( A => v_KEY32_IN_1_port, B => n162, C => n8279, D => 
                           v_TEMP_VECTOR_1_port, Z => n218);
   U799 : AO3 port map( A => n208, B => n159, C => n209, D => n210, Z => n6693)
                           ;
   U800 : AO2 port map( A => v_KEY32_IN_2_port, B => n162, C => n8279, D => 
                           v_TEMP_VECTOR_2_port, Z => n210);
   U801 : AO3 port map( A => n159, B => n199, C => n200, D => n201, Z => n6692)
                           ;
   U802 : AO2 port map( A => v_KEY32_IN_3_port, B => n162, C => n8279, D => 
                           v_TEMP_VECTOR_3_port, Z => n201);
   U803 : AO3 port map( A => n159, B => n191, C => n192, D => n193, Z => n6691)
                           ;
   U804 : AO2 port map( A => v_KEY32_IN_4_port, B => n162, C => n8279, D => 
                           v_TEMP_VECTOR_4_port, Z => n193);
   U805 : AO3 port map( A => n183, B => n159, C => n184, D => n185, Z => n6690)
                           ;
   U806 : AO2 port map( A => v_KEY32_IN_5_port, B => n162, C => n8279, D => 
                           v_TEMP_VECTOR_5_port, Z => n185);
   U807 : AO7 port map( A => n2004, B => n172, C => n173, Z => n6689);
   U808 : AO2 port map( A => n2297, B => n174, C => v_KEY32_IN_6_port, D => 
                           n162, Z => n173);
   U809 : AO3 port map( A => n158, B => n159, C => n160, D => n161, Z => n6688)
                           ;
   U810 : AO2 port map( A => v_KEY32_IN_7_port, B => n162, C => n8279, D => 
                           v_TEMP_VECTOR_7_port, Z => n161);
   U811 : AO7 port map( A => v_KEY_COL_OUT0_8_port, B => n2300, C => n8275, Z 
                           => n152);
   U812 : AO7 port map( A => v_KEY_COL_OUT0_16_port, B => n2302, C => n8277, Z 
                           => n111);
   U813 : AO7 port map( A => v_KEY_COL_OUT0_24_port, B => n2304, C => n8220, Z 
                           => n61);
   U814 : AO7 port map( A => v_KEY_COL_OUT0_9_port, B => n2300, C => n8275, Z 
                           => n146);
   U815 : AO7 port map( A => v_KEY_COL_OUT0_17_port, B => n2302, C => n8277, Z 
                           => n105);
   U816 : AO7 port map( A => v_KEY_COL_OUT0_25_port, B => n2304, C => n8220, Z 
                           => n52);
   U817 : AO7 port map( A => v_KEY_COL_OUT0_10_port, B => n2299, C => n8275, Z 
                           => n142);
   U818 : AO7 port map( A => v_KEY_COL_OUT0_18_port, B => n2301, C => n8277, Z 
                           => n101);
   U819 : AO7 port map( A => v_KEY_COL_OUT0_26_port, B => n2303, C => n8220, Z 
                           => n47);
   U820 : AO7 port map( A => v_KEY_COL_OUT0_11_port, B => n2299, C => n8275, Z 
                           => n138);
   U821 : AO7 port map( A => v_KEY_COL_OUT0_19_port, B => n2301, C => n8277, Z 
                           => n97);
   U823 : AO7 port map( A => v_KEY_COL_OUT0_27_port, B => n2303, C => n8220, Z 
                           => n42);
   U824 : AO7 port map( A => v_KEY_COL_OUT0_12_port, B => n2299, C => n8275, Z 
                           => n134);
   U825 : AO7 port map( A => v_KEY_COL_OUT0_20_port, B => n2301, C => n8277, Z 
                           => n93);
   U826 : AO7 port map( A => v_KEY_COL_OUT0_28_port, B => n2303, C => n8220, Z 
                           => n37);
   U827 : AO7 port map( A => v_KEY_COL_OUT0_13_port, B => n2299, C => n8275, Z 
                           => n130);
   U828 : AO7 port map( A => v_KEY_COL_OUT0_21_port, B => n2301, C => n8277, Z 
                           => n89);
   U829 : AO7 port map( A => v_KEY_COL_OUT0_29_port, B => n2303, C => n8220, Z 
                           => n32);
   U830 : AO7 port map( A => v_KEY_COL_OUT0_14_port, B => n2299, C => n8275, Z 
                           => n126);
   U831 : AO7 port map( A => v_KEY_COL_OUT0_22_port, B => n2301, C => n8277, Z 
                           => n85);
   U832 : AO7 port map( A => v_KEY_COL_OUT0_30_port, B => n2303, C => n8220, Z 
                           => n27);
   U833 : AO7 port map( A => v_KEY_COL_OUT0_15_port, B => n2299, C => n8275, Z 
                           => n120);
   U834 : AO7 port map( A => v_KEY_COL_OUT0_23_port, B => n2301, C => n8277, Z 
                           => n79);
   U835 : AO7 port map( A => v_KEY_COL_OUT0_31_port, B => n2303, C => n8220, Z 
                           => n20);
   U836 : AO3 port map( A => n1954, B => n114, C => n147, D => n148, Z => n6687
                           );
   U837 : AO2 port map( A => n151, B => v_KEY_COL_OUT0_8_port, C => 
                           v_TEMP_VECTOR_8_port, D => n152, Z => n147);
   U838 : AO2 port map( A => n117, B => v_TEMP_VECTOR_16_port, C => 
                           v_KEY32_IN_8_port, D => n118, Z => n148);
   U839 : AO3 port map( A => n1954, B => n73, C => n106, D => n107, Z => n6679)
                           ;
   U840 : AO2 port map( A => n110, B => v_KEY_COL_OUT0_16_port, C => 
                           v_TEMP_VECTOR_16_port, D => n111, Z => n106);
   U841 : AO2 port map( A => n76, B => v_TEMP_VECTOR_24_port, C => 
                           v_KEY32_IN_16_port, D => n77, Z => n107);
   U842 : AO3 port map( A => n13, B => n1954, C => n54, D => n55, Z => n6671);
   U843 : AO2 port map( A => n60, B => v_KEY_COL_OUT0_24_port, C => 
                           v_TEMP_VECTOR_24_port, D => n61, Z => n54);
   U844 : AO2 port map( A => v_TEMP_VECTOR_0_port, B => n17, C => 
                           v_KEY32_IN_24_port, D => n18, Z => n55);
   U845 : AO3 port map( A => n1955, B => n114, C => n143, D => n144, Z => n6686
                           );
   U846 : AO2 port map( A => n145, B => v_KEY_COL_OUT0_9_port, C => 
                           v_TEMP_VECTOR_9_port, D => n146, Z => n143);
   U847 : AO2 port map( A => n117, B => v_TEMP_VECTOR_17_port, C => 
                           v_KEY32_IN_9_port, D => n118, Z => n144);
   U848 : AO3 port map( A => n1955, B => n73, C => n102, D => n103, Z => n6678)
                           ;
   U849 : AO2 port map( A => n104, B => v_KEY_COL_OUT0_17_port, C => 
                           v_TEMP_VECTOR_17_port, D => n105, Z => n102);
   U850 : AO2 port map( A => n76, B => v_TEMP_VECTOR_25_port, C => 
                           v_KEY32_IN_17_port, D => n77, Z => n103);
   U851 : AO3 port map( A => n13, B => n1955, C => n49, D => n50, Z => n6670);
   U852 : AO2 port map( A => n51, B => v_KEY_COL_OUT0_25_port, C => 
                           v_TEMP_VECTOR_25_port, D => n52, Z => n49);
   U853 : AO2 port map( A => v_TEMP_VECTOR_1_port, B => n17, C => 
                           v_KEY32_IN_25_port, D => n18, Z => n50);
   U854 : AO3 port map( A => n1978, B => n114, C => n139, D => n140, Z => n6685
                           );
   U855 : AO2 port map( A => n141, B => v_KEY_COL_OUT0_10_port, C => 
                           v_TEMP_VECTOR_10_port, D => n142, Z => n139);
   U856 : AO2 port map( A => n117, B => v_TEMP_VECTOR_18_port, C => 
                           v_KEY32_IN_10_port, D => n118, Z => n140);
   U857 : AO3 port map( A => n1978, B => n73, C => n98, D => n99, Z => n6677);
   U858 : AO2 port map( A => n100, B => v_KEY_COL_OUT0_18_port, C => 
                           v_TEMP_VECTOR_18_port, D => n101, Z => n98);
   U859 : AO2 port map( A => n76, B => v_TEMP_VECTOR_26_port, C => 
                           v_KEY32_IN_18_port, D => n77, Z => n99);
   U860 : AO3 port map( A => n13, B => n1978, C => n44, D => n45, Z => n6669);
   U861 : AO2 port map( A => n46, B => v_KEY_COL_OUT0_26_port, C => 
                           v_TEMP_VECTOR_26_port, D => n47, Z => n44);
   U862 : AO2 port map( A => v_TEMP_VECTOR_2_port, B => n17, C => 
                           v_KEY32_IN_26_port, D => n18, Z => n45);
   U863 : AO3 port map( A => n1976, B => n114, C => n135, D => n136, Z => n6684
                           );
   U864 : AO2 port map( A => n137, B => v_KEY_COL_OUT0_11_port, C => 
                           v_TEMP_VECTOR_11_port, D => n138, Z => n135);
   U865 : AO2 port map( A => n117, B => v_TEMP_VECTOR_19_port, C => 
                           v_KEY32_IN_11_port, D => n118, Z => n136);
   U867 : AO3 port map( A => n1976, B => n73, C => n94, D => n95, Z => n6676);
   U868 : AO2 port map( A => n96, B => v_KEY_COL_OUT0_19_port, C => 
                           v_TEMP_VECTOR_19_port, D => n97, Z => n94);
   U869 : AO2 port map( A => n76, B => v_TEMP_VECTOR_27_port, C => 
                           v_KEY32_IN_19_port, D => n77, Z => n95);
   U870 : AO3 port map( A => n13, B => n1976, C => n39, D => n40, Z => n6668);
   U871 : AO2 port map( A => n41, B => v_KEY_COL_OUT0_27_port, C => 
                           v_TEMP_VECTOR_27_port, D => n42, Z => n39);
   U872 : AO2 port map( A => v_TEMP_VECTOR_3_port, B => n17, C => 
                           v_KEY32_IN_27_port, D => n18, Z => n40);
   U873 : AO3 port map( A => n1974, B => n114, C => n131, D => n132, Z => n6683
                           );
   U874 : AO2 port map( A => n133, B => v_KEY_COL_OUT0_12_port, C => 
                           v_TEMP_VECTOR_12_port, D => n134, Z => n131);
   U875 : AO2 port map( A => n117, B => v_TEMP_VECTOR_20_port, C => 
                           v_KEY32_IN_12_port, D => n118, Z => n132);
   U876 : AO3 port map( A => n1974, B => n73, C => n90, D => n91, Z => n6675);
   U877 : AO2 port map( A => n92, B => v_KEY_COL_OUT0_20_port, C => 
                           v_TEMP_VECTOR_20_port, D => n93, Z => n90);
   U878 : AO2 port map( A => n76, B => v_TEMP_VECTOR_28_port, C => 
                           v_KEY32_IN_20_port, D => n77, Z => n91);
   U879 : AO3 port map( A => n13, B => n1974, C => n34, D => n35, Z => n6667);
   U880 : AO2 port map( A => n36, B => v_KEY_COL_OUT0_28_port, C => 
                           v_TEMP_VECTOR_28_port, D => n37, Z => n34);
   U881 : AO2 port map( A => v_TEMP_VECTOR_4_port, B => n17, C => 
                           v_KEY32_IN_28_port, D => n18, Z => n35);
   U882 : AO3 port map( A => n1964, B => n114, C => n127, D => n128, Z => n6682
                           );
   U883 : AO2 port map( A => n129, B => v_KEY_COL_OUT0_13_port, C => 
                           v_TEMP_VECTOR_13_port, D => n130, Z => n127);
   U884 : AO2 port map( A => n117, B => v_TEMP_VECTOR_21_port, C => 
                           v_KEY32_IN_13_port, D => n118, Z => n128);
   U885 : AO3 port map( A => n1964, B => n73, C => n86, D => n87, Z => n6674);
   U886 : AO2 port map( A => n88, B => v_KEY_COL_OUT0_21_port, C => 
                           v_TEMP_VECTOR_21_port, D => n89, Z => n86);
   U887 : AO2 port map( A => n76, B => v_TEMP_VECTOR_29_port, C => 
                           v_KEY32_IN_21_port, D => n77, Z => n87);
   U888 : AO3 port map( A => n13, B => n1964, C => n29, D => n30, Z => n6666);
   U889 : AO2 port map( A => n31, B => v_KEY_COL_OUT0_29_port, C => 
                           v_TEMP_VECTOR_29_port, D => n32, Z => n29);
   U890 : AO2 port map( A => v_TEMP_VECTOR_5_port, B => n17, C => 
                           v_KEY32_IN_29_port, D => n18, Z => n30);
   U891 : AO3 port map( A => n1959, B => n114, C => n123, D => n124, Z => n6681
                           );
   U892 : AO2 port map( A => n125, B => v_KEY_COL_OUT0_14_port, C => 
                           v_TEMP_VECTOR_14_port, D => n126, Z => n123);
   U893 : AO2 port map( A => n117, B => v_TEMP_VECTOR_22_port, C => 
                           v_KEY32_IN_14_port, D => n118, Z => n124);
   U894 : AO3 port map( A => n1959, B => n73, C => n82, D => n83, Z => n6673);
   U895 : AO2 port map( A => n84, B => v_KEY_COL_OUT0_22_port, C => 
                           v_TEMP_VECTOR_22_port, D => n85, Z => n82);
   U896 : AO2 port map( A => n76, B => v_TEMP_VECTOR_30_port, C => 
                           v_KEY32_IN_22_port, D => n77, Z => n83);
   U897 : AO3 port map( A => n13, B => n1959, C => n24, D => n25, Z => n6665);
   U898 : AO2 port map( A => n26, B => v_KEY_COL_OUT0_30_port, C => 
                           v_TEMP_VECTOR_30_port, D => n27, Z => n24);
   U899 : AO2 port map( A => v_TEMP_VECTOR_6_port, B => n17, C => 
                           v_KEY32_IN_30_port, D => n18, Z => n25);
   U900 : AO3 port map( A => n1960, B => n114, C => n115, D => n116, Z => n6680
                           );
   U901 : AO2 port map( A => n119, B => v_KEY_COL_OUT0_15_port, C => 
                           v_TEMP_VECTOR_15_port, D => n120, Z => n115);
   U902 : AO2 port map( A => n117, B => v_TEMP_VECTOR_23_port, C => 
                           v_KEY32_IN_15_port, D => n118, Z => n116);
   U903 : AO3 port map( A => n1960, B => n73, C => n74, D => n75, Z => n6672);
   U904 : AO2 port map( A => n78, B => v_KEY_COL_OUT0_23_port, C => 
                           v_TEMP_VECTOR_23_port, D => n79, Z => n74);
   U905 : AO2 port map( A => n76, B => v_TEMP_VECTOR_31_port, C => 
                           v_KEY32_IN_23_port, D => n77, Z => n75);
   U906 : AO3 port map( A => n13, B => n1960, C => n15, D => n16, Z => n6664);
   U907 : AO2 port map( A => n19, B => v_KEY_COL_OUT0_31_port, C => 
                           v_TEMP_VECTOR_31_port, D => n20, Z => n15);
   U908 : AO2 port map( A => v_TEMP_VECTOR_7_port, B => n17, C => 
                           v_KEY32_IN_31_port, D => n18, Z => n16);
   U909 : AO2 port map( A => v_TEMP_VECTOR_30_port, B => n2166, C => 
                           v_TEMP_VECTOR_22_port, D => n2168, Z => n2246);
   U911 : IVDA port map( A => n1997, Y => n381, Z => n2214);
   U912 : AO2 port map( A => v_TEMP_VECTOR_24_port, B => n2166, C => 
                           v_TEMP_VECTOR_16_port, D => n2168, Z => n2265);
   U913 : AO2 port map( A => v_KEY32_IN_8_port, B => n266, C => 
                           v_TEMP_VECTOR_8_port, D => n271, Z => n2428);
   U914 : AO2 port map( A => v_KEY32_IN_16_port, B => n266, C => 
                           v_TEMP_VECTOR_16_port, D => n271, Z => n2436);
   U915 : AO2 port map( A => v_KEY32_IN_24_port, B => n266, C => 
                           v_TEMP_VECTOR_24_port, D => n271, Z => n2444);
   U916 : AO2 port map( A => v_KEY32_IN_9_port, B => n266, C => 
                           v_TEMP_VECTOR_9_port, D => n271, Z => n2429);
   U917 : AO2 port map( A => v_KEY32_IN_17_port, B => n266, C => 
                           v_TEMP_VECTOR_17_port, D => n271, Z => n2437);
   U918 : AO2 port map( A => v_KEY32_IN_25_port, B => n266, C => 
                           v_TEMP_VECTOR_25_port, D => n271, Z => n2445);
   U919 : AO2 port map( A => v_KEY32_IN_10_port, B => n266, C => 
                           v_TEMP_VECTOR_10_port, D => n271, Z => n2430);
   U920 : AO2 port map( A => v_KEY32_IN_18_port, B => n266, C => 
                           v_TEMP_VECTOR_18_port, D => n271, Z => n2438);
   U921 : AO2 port map( A => v_KEY32_IN_26_port, B => n266, C => 
                           v_TEMP_VECTOR_26_port, D => n271, Z => n2446);
   U922 : AO2 port map( A => v_KEY32_IN_11_port, B => n266, C => 
                           v_TEMP_VECTOR_11_port, D => n271, Z => n2431);
   U923 : AO2 port map( A => v_KEY32_IN_19_port, B => n266, C => 
                           v_TEMP_VECTOR_19_port, D => n271, Z => n2439);
   U924 : AO2 port map( A => v_KEY32_IN_27_port, B => n266, C => 
                           v_TEMP_VECTOR_27_port, D => n271, Z => n2447);
   U925 : AO2 port map( A => v_KEY32_IN_12_port, B => n266, C => 
                           v_TEMP_VECTOR_12_port, D => n271, Z => n2432);
   U926 : AO2 port map( A => v_KEY32_IN_20_port, B => n266, C => 
                           v_TEMP_VECTOR_20_port, D => n271, Z => n2440);
   U927 : AO2 port map( A => v_KEY32_IN_28_port, B => n266, C => 
                           v_TEMP_VECTOR_28_port, D => n271, Z => n2448);
   U928 : AO2 port map( A => v_KEY32_IN_4_port, B => n266, C => 
                           v_TEMP_VECTOR_4_port, D => n271, Z => n2424);
   U929 : AO2 port map( A => v_KEY32_IN_13_port, B => n266, C => 
                           v_TEMP_VECTOR_13_port, D => n271, Z => n2433);
   U930 : AO2 port map( A => v_KEY32_IN_21_port, B => n266, C => 
                           v_TEMP_VECTOR_21_port, D => n271, Z => n2441);
   U931 : AO2 port map( A => v_KEY32_IN_29_port, B => n266, C => 
                           v_TEMP_VECTOR_29_port, D => n271, Z => n2449);
   U932 : AO2 port map( A => v_KEY32_IN_5_port, B => n266, C => 
                           v_TEMP_VECTOR_5_port, D => n271, Z => n2425);
   U933 : AO2 port map( A => v_KEY32_IN_14_port, B => n266, C => 
                           v_TEMP_VECTOR_14_port, D => n271, Z => n2434);
   U934 : AO2 port map( A => v_KEY32_IN_22_port, B => n266, C => 
                           v_TEMP_VECTOR_22_port, D => n271, Z => n2442);
   U935 : AO2 port map( A => v_KEY32_IN_30_port, B => n266, C => 
                           v_TEMP_VECTOR_30_port, D => n271, Z => n2450);
   U936 : AO2 port map( A => v_KEY32_IN_6_port, B => n266, C => 
                           v_TEMP_VECTOR_6_port, D => n271, Z => n2426);
   U937 : AO2 port map( A => v_KEY32_IN_15_port, B => n266, C => 
                           v_TEMP_VECTOR_15_port, D => n271, Z => n2435);
   U938 : AO2 port map( A => v_KEY32_IN_23_port, B => n266, C => 
                           v_TEMP_VECTOR_23_port, D => n271, Z => n2443);
   U939 : AO2 port map( A => v_KEY32_IN_31_port, B => n266, C => 
                           v_TEMP_VECTOR_31_port, D => n271, Z => n2451);
   U940 : AO2 port map( A => v_KEY32_IN_7_port, B => n266, C => 
                           v_TEMP_VECTOR_7_port, D => n271, Z => n2427);
   U941 : AO4 port map( A => n2530, B => n8054, C => n6731, D => n8048, Z => 
                           n5102);
   U942 : AO4 port map( A => n2531, B => n8034, C => n6731, D => n8028, Z => 
                           n5103);
   U943 : AO4 port map( A => n2528, B => n8014, C => n6731, D => n8008, Z => 
                           n5104);
   U944 : AO4 port map( A => n2529, B => n7994, C => n6731, D => n7988, Z => 
                           n5105);
   U945 : AO4 port map( A => n2526, B => n7974, C => n6731, D => n7968, Z => 
                           n5106);
   U946 : AO4 port map( A => n2527, B => n7954, C => n6731, D => n7948, Z => 
                           n5107);
   U947 : AO4 port map( A => n2524, B => n7934, C => n6731, D => n7928, Z => 
                           n5108);
   U948 : AO4 port map( A => n2525, B => n7914, C => n6731, D => n7908, Z => 
                           n5109);
   U949 : AO4 port map( A => n2594, B => n8055, C => n2401, D => n8044, Z => 
                           n5614);
   U950 : AO4 port map( A => n2595, B => n8035, C => n2401, D => n8024, Z => 
                           n5615);
   U951 : AO4 port map( A => n2592, B => n8015, C => n2401, D => n8004, Z => 
                           n5616);
   U952 : AO4 port map( A => n2593, B => n7995, C => n2401, D => n7984, Z => 
                           n5617);
   U953 : AO4 port map( A => n2590, B => n7975, C => n2401, D => n7964, Z => 
                           n5618);
   U955 : AO4 port map( A => n2591, B => n7955, C => n2401, D => n7944, Z => 
                           n5619);
   U956 : AO4 port map( A => n2588, B => n7935, C => n2401, D => n7924, Z => 
                           n5620);
   U957 : AO4 port map( A => n2589, B => n7915, C => n2401, D => n7904, Z => 
                           n5621);
   U958 : AO4 port map( A => n2658, B => n8055, C => n2353, D => n8040, Z => 
                           n6126);
   U959 : AO4 port map( A => n2659, B => n8035, C => n2353, D => n8020, Z => 
                           n6127);
   U960 : AO4 port map( A => n2656, B => n8015, C => n2353, D => n8000, Z => 
                           n6128);
   U961 : AO4 port map( A => n2657, B => n7995, C => n2353, D => n7980, Z => 
                           n6129);
   U962 : AO4 port map( A => n2654, B => n7975, C => n2353, D => n7960, Z => 
                           n6130);
   U963 : AO4 port map( A => n2655, B => n7955, C => n2353, D => n7940, Z => 
                           n6131);
   U964 : AO4 port map( A => n2652, B => n7935, C => n2353, D => n7920, Z => 
                           n6132);
   U965 : AO4 port map( A => n2653, B => n7915, C => n2353, D => n7900, Z => 
                           n6133);
   U966 : AO4 port map( A => n2787, B => n8054, C => n6725, D => n8048, Z => 
                           n5166);
   U967 : AO4 port map( A => n2788, B => n8034, C => n6725, D => n8028, Z => 
                           n5167);
   U968 : AO4 port map( A => n2785, B => n8014, C => n6725, D => n8008, Z => 
                           n5168);
   U969 : AO4 port map( A => n2786, B => n7994, C => n6725, D => n7988, Z => 
                           n5169);
   U970 : AO4 port map( A => n2783, B => n7974, C => n6725, D => n7968, Z => 
                           n5170);
   U971 : AO4 port map( A => n2784, B => n7954, C => n6725, D => n7948, Z => 
                           n5171);
   U972 : AO4 port map( A => n2781, B => n7934, C => n6725, D => n7928, Z => 
                           n5172);
   U973 : AO4 port map( A => n2782, B => n7914, C => n6725, D => n7908, Z => 
                           n5173);
   U974 : AO4 port map( A => n2851, B => n8055, C => n2395, D => n8044, Z => 
                           n5678);
   U975 : AO4 port map( A => n2852, B => n8035, C => n2395, D => n8024, Z => 
                           n5679);
   U976 : AO4 port map( A => n2849, B => n8015, C => n2395, D => n8004, Z => 
                           n5680);
   U977 : AO4 port map( A => n2850, B => n7995, C => n2395, D => n7984, Z => 
                           n5681);
   U978 : AO4 port map( A => n2847, B => n7975, C => n2395, D => n7964, Z => 
                           n5682);
   U979 : AO4 port map( A => n2848, B => n7955, C => n2395, D => n7944, Z => 
                           n5683);
   U980 : AO4 port map( A => n2845, B => n7935, C => n2395, D => n7924, Z => 
                           n5684);
   U981 : AO4 port map( A => n2846, B => n7915, C => n2395, D => n7904, Z => 
                           n5685);
   U982 : AO4 port map( A => n2915, B => n8055, C => n2347, D => n8040, Z => 
                           n6190);
   U983 : AO4 port map( A => n2916, B => n8035, C => n2347, D => n8020, Z => 
                           n6191);
   U984 : AO4 port map( A => n2913, B => n8015, C => n2347, D => n8000, Z => 
                           n6192);
   U985 : AO4 port map( A => n2914, B => n7995, C => n2347, D => n7980, Z => 
                           n6193);
   U986 : AO4 port map( A => n2911, B => n7975, C => n2347, D => n7960, Z => 
                           n6194);
   U987 : AO4 port map( A => n2912, B => n7955, C => n2347, D => n7940, Z => 
                           n6195);
   U988 : AO4 port map( A => n2909, B => n7935, C => n2347, D => n7920, Z => 
                           n6196);
   U989 : AO4 port map( A => n2910, B => n7915, C => n2347, D => n7900, Z => 
                           n6197);
   U990 : AO4 port map( A => n3043, B => n8054, C => n6719, D => n8047, Z => 
                           n5230);
   U991 : AO4 port map( A => n3044, B => n8034, C => n6719, D => n8027, Z => 
                           n5231);
   U992 : AO4 port map( A => n3041, B => n8014, C => n6719, D => n8007, Z => 
                           n5232);
   U993 : AO4 port map( A => n3042, B => n7994, C => n6719, D => n7987, Z => 
                           n5233);
   U994 : AO4 port map( A => n3039, B => n7974, C => n6719, D => n7967, Z => 
                           n5234);
   U995 : AO4 port map( A => n3040, B => n7954, C => n6719, D => n7947, Z => 
                           n5235);
   U996 : AO4 port map( A => n3037, B => n7934, C => n6719, D => n7927, Z => 
                           n5236);
   U997 : AO4 port map( A => n3038, B => n7914, C => n6719, D => n7907, Z => 
                           n5237);
   U999 : AO4 port map( A => n3107, B => n8055, C => n2389, D => n8043, Z => 
                           n5742);
   U1000 : AO4 port map( A => n3108, B => n8035, C => n2389, D => n8023, Z => 
                           n5743);
   U1001 : AO4 port map( A => n3105, B => n8015, C => n2389, D => n8003, Z => 
                           n5744);
   U1002 : AO4 port map( A => n3106, B => n7995, C => n2389, D => n7983, Z => 
                           n5745);
   U1003 : AO4 port map( A => n3103, B => n7975, C => n2389, D => n7963, Z => 
                           n5746);
   U1004 : AO4 port map( A => n3104, B => n7955, C => n2389, D => n7943, Z => 
                           n5747);
   U1005 : AO4 port map( A => n3101, B => n7935, C => n2389, D => n7923, Z => 
                           n5748);
   U1006 : AO4 port map( A => n3102, B => n7915, C => n2389, D => n7903, Z => 
                           n5749);
   U1007 : AO4 port map( A => n3171, B => n8055, C => n2341, D => n8039, Z => 
                           n6254);
   U1008 : AO4 port map( A => n3172, B => n8035, C => n2341, D => n8019, Z => 
                           n6255);
   U1009 : AO4 port map( A => n3169, B => n8015, C => n2341, D => n7999, Z => 
                           n6256);
   U1010 : AO4 port map( A => n3170, B => n7995, C => n2341, D => n7979, Z => 
                           n6257);
   U1011 : AO4 port map( A => n3167, B => n7975, C => n2341, D => n7959, Z => 
                           n6258);
   U1012 : AO4 port map( A => n3168, B => n7955, C => n2341, D => n7939, Z => 
                           n6259);
   U1013 : AO4 port map( A => n3165, B => n7935, C => n2341, D => n7919, Z => 
                           n6260);
   U1014 : AO4 port map( A => n3166, B => n7915, C => n2341, D => n7899, Z => 
                           n6261);
   U1015 : AO4 port map( A => n3299, B => n8054, C => n6656, D => n8047, Z => 
                           n5294);
   U1016 : AO4 port map( A => n3300, B => n8034, C => n6656, D => n8027, Z => 
                           n5295);
   U1017 : AO4 port map( A => n3297, B => n8014, C => n6656, D => n8007, Z => 
                           n5296);
   U1018 : AO4 port map( A => n3298, B => n7994, C => n6656, D => n7987, Z => 
                           n5297);
   U1019 : AO4 port map( A => n3295, B => n7974, C => n6656, D => n7967, Z => 
                           n5298);
   U1020 : AO4 port map( A => n3296, B => n7954, C => n6656, D => n7947, Z => 
                           n5299);
   U1021 : AO4 port map( A => n3293, B => n7934, C => n6656, D => n7927, Z => 
                           n5300);
   U1022 : AO4 port map( A => n3294, B => n7914, C => n6656, D => n7907, Z => 
                           n5301);
   U1023 : AO4 port map( A => n3363, B => n8055, C => n2383, D => n8043, Z => 
                           n5806);
   U1024 : AO4 port map( A => n3364, B => n8035, C => n2383, D => n8023, Z => 
                           n5807);
   U1025 : AO4 port map( A => n3361, B => n8015, C => n2383, D => n8003, Z => 
                           n5808);
   U1026 : AO4 port map( A => n3362, B => n7995, C => n2383, D => n7983, Z => 
                           n5809);
   U1027 : AO4 port map( A => n3359, B => n7975, C => n2383, D => n7963, Z => 
                           n5810);
   U1028 : AO4 port map( A => n3360, B => n7955, C => n2383, D => n7943, Z => 
                           n5811);
   U1029 : AO4 port map( A => n3357, B => n7935, C => n2383, D => n7923, Z => 
                           n5812);
   U1030 : AO4 port map( A => n3358, B => n7915, C => n2383, D => n7903, Z => 
                           n5813);
   U1031 : AO4 port map( A => n3427, B => n8055, C => n2335, D => n8039, Z => 
                           n6318);
   U1032 : AO4 port map( A => n3428, B => n8035, C => n2335, D => n8019, Z => 
                           n6319);
   U1033 : AO4 port map( A => n3425, B => n8015, C => n2335, D => n7999, Z => 
                           n6320);
   U1034 : AO4 port map( A => n3426, B => n7995, C => n2335, D => n7979, Z => 
                           n6321);
   U1035 : AO4 port map( A => n3423, B => n7975, C => n2335, D => n7959, Z => 
                           n6322);
   U1036 : AO4 port map( A => n3424, B => n7955, C => n2335, D => n7939, Z => 
                           n6323);
   U1037 : AO4 port map( A => n3421, B => n7935, C => n2335, D => n7919, Z => 
                           n6324);
   U1038 : AO4 port map( A => n3422, B => n7915, C => n2335, D => n7899, Z => 
                           n6325);
   U1039 : AO4 port map( A => n3555, B => n8054, C => n2480, D => n8046, Z => 
                           n5358);
   U1040 : AO4 port map( A => n3556, B => n8034, C => n2480, D => n8026, Z => 
                           n5359);
   U1041 : AO4 port map( A => n3553, B => n8014, C => n2480, D => n8006, Z => 
                           n5360);
   U1043 : AO4 port map( A => n3554, B => n7994, C => n2480, D => n7986, Z => 
                           n5361);
   U1044 : AO4 port map( A => n3551, B => n7974, C => n2480, D => n7966, Z => 
                           n5362);
   U1045 : AO4 port map( A => n3552, B => n7954, C => n2480, D => n7946, Z => 
                           n5363);
   U1046 : AO4 port map( A => n3549, B => n7934, C => n2480, D => n7926, Z => 
                           n5364);
   U1047 : AO4 port map( A => n3550, B => n7914, C => n2480, D => n7906, Z => 
                           n5365);
   U1048 : AO4 port map( A => n3619, B => n8055, C => n2377, D => n8042, Z => 
                           n5870);
   U1049 : AO4 port map( A => n3620, B => n8035, C => n2377, D => n8022, Z => 
                           n5871);
   U1050 : AO4 port map( A => n3617, B => n8015, C => n2377, D => n8002, Z => 
                           n5872);
   U1051 : AO4 port map( A => n3618, B => n7995, C => n2377, D => n7982, Z => 
                           n5873);
   U1052 : AO4 port map( A => n3615, B => n7975, C => n2377, D => n7962, Z => 
                           n5874);
   U1053 : AO4 port map( A => n3616, B => n7955, C => n2377, D => n7942, Z => 
                           n5875);
   U1054 : AO4 port map( A => n3613, B => n7935, C => n2377, D => n7922, Z => 
                           n5876);
   U1055 : AO4 port map( A => n3614, B => n7915, C => n2377, D => n7902, Z => 
                           n5877);
   U1056 : AO4 port map( A => n3683, B => n8056, C => n2329, D => n8038, Z => 
                           n6382);
   U1057 : AO4 port map( A => n3684, B => n8036, C => n2329, D => n8018, Z => 
                           n6383);
   U1058 : AO4 port map( A => n3681, B => n8016, C => n2329, D => n7998, Z => 
                           n6384);
   U1059 : AO4 port map( A => n3682, B => n7996, C => n2329, D => n7978, Z => 
                           n6385);
   U1060 : AO4 port map( A => n3679, B => n7976, C => n2329, D => n7958, Z => 
                           n6386);
   U1061 : AO4 port map( A => n3680, B => n7956, C => n2329, D => n7938, Z => 
                           n6387);
   U1062 : AO4 port map( A => n3677, B => n7936, C => n2329, D => n7918, Z => 
                           n6388);
   U1063 : AO4 port map( A => n3678, B => n7916, C => n2329, D => n7898, Z => 
                           n6389);
   U1064 : AO4 port map( A => n3747, B => n8054, C => n6757, D => n8050, Z => 
                           n4846);
   U1065 : AO4 port map( A => n3748, B => n8034, C => n6757, D => n8030, Z => 
                           n4847);
   U1066 : AO4 port map( A => n3745, B => n8014, C => n6757, D => n8010, Z => 
                           n4848);
   U1067 : AO4 port map( A => n3746, B => n7994, C => n6757, D => n7990, Z => 
                           n4849);
   U1068 : AO4 port map( A => n3743, B => n7974, C => n6757, D => n7970, Z => 
                           n4850);
   U1069 : AO4 port map( A => n3744, B => n7954, C => n6757, D => n7950, Z => 
                           n4851);
   U1070 : AO4 port map( A => n3741, B => n7934, C => n6757, D => n7930, Z => 
                           n4852);
   U1071 : AO4 port map( A => n3742, B => n7914, C => n6757, D => n7910, Z => 
                           n4853);
   U1072 : AO4 port map( A => n3811, B => n8054, C => n2419, D => n8046, Z => 
                           n5422);
   U1073 : AO4 port map( A => n3812, B => n8034, C => n2419, D => n8026, Z => 
                           n5423);
   U1074 : AO4 port map( A => n3809, B => n8014, C => n2419, D => n8006, Z => 
                           n5424);
   U1075 : AO4 port map( A => n3810, B => n7994, C => n2419, D => n7986, Z => 
                           n5425);
   U1076 : AO4 port map( A => n3807, B => n7974, C => n2419, D => n7966, Z => 
                           n5426);
   U1077 : AO4 port map( A => n3808, B => n7954, C => n2419, D => n7946, Z => 
                           n5427);
   U1078 : AO4 port map( A => n3805, B => n7934, C => n2419, D => n7926, Z => 
                           n5428);
   U1079 : AO4 port map( A => n3806, B => n7914, C => n2419, D => n7906, Z => 
                           n5429);
   U1080 : AO4 port map( A => n3875, B => n8055, C => n2371, D => n8042, Z => 
                           n5934);
   U1081 : AO4 port map( A => n3876, B => n8035, C => n2371, D => n8022, Z => 
                           n5935);
   U1082 : AO4 port map( A => n3873, B => n8015, C => n2371, D => n8002, Z => 
                           n5936);
   U1083 : AO4 port map( A => n3874, B => n7995, C => n2371, D => n7982, Z => 
                           n5937);
   U1084 : AO4 port map( A => n3871, B => n7975, C => n2371, D => n7962, Z => 
                           n5938);
   U1085 : AO4 port map( A => n3872, B => n7955, C => n2371, D => n7942, Z => 
                           n5939);
   U1087 : AO4 port map( A => n3869, B => n7935, C => n2371, D => n7922, Z => 
                           n5940);
   U1088 : AO4 port map( A => n3870, B => n7915, C => n2371, D => n7902, Z => 
                           n5941);
   U1089 : AO4 port map( A => n3939, B => n8056, C => n2323, D => n8038, Z => 
                           n6446);
   U1090 : AO4 port map( A => n3940, B => n8036, C => n2323, D => n8018, Z => 
                           n6447);
   U1091 : AO4 port map( A => n3937, B => n8016, C => n2323, D => n7998, Z => 
                           n6448);
   U1092 : AO4 port map( A => n3938, B => n7996, C => n2323, D => n7978, Z => 
                           n6449);
   U1093 : AO4 port map( A => n3935, B => n7976, C => n2323, D => n7958, Z => 
                           n6450);
   U1094 : AO4 port map( A => n3936, B => n7956, C => n2323, D => n7938, Z => 
                           n6451);
   U1095 : AO4 port map( A => n3933, B => n7936, C => n2323, D => n7918, Z => 
                           n6452);
   U1096 : AO4 port map( A => n3934, B => n7916, C => n2323, D => n7898, Z => 
                           n6453);
   U1097 : AO4 port map( A => n4003, B => n8054, C => n6751, D => n8050, Z => 
                           n4910);
   U1098 : AO4 port map( A => n4004, B => n8034, C => n6751, D => n8030, Z => 
                           n4911);
   U1099 : AO4 port map( A => n4001, B => n8014, C => n6751, D => n8010, Z => 
                           n4912);
   U1100 : AO4 port map( A => n4002, B => n7994, C => n6751, D => n7990, Z => 
                           n4913);
   U1101 : AO4 port map( A => n3999, B => n7974, C => n6751, D => n7970, Z => 
                           n4914);
   U1102 : AO4 port map( A => n4000, B => n7954, C => n6751, D => n7950, Z => 
                           n4915);
   U1103 : AO4 port map( A => n3997, B => n7934, C => n6751, D => n7930, Z => 
                           n4916);
   U1104 : AO4 port map( A => n3998, B => n7914, C => n6751, D => n7910, Z => 
                           n4917);
   U1105 : AO4 port map( A => n4067, B => n8055, C => n2413, D => n8045, Z => 
                           n5486);
   U1106 : AO4 port map( A => n4068, B => n8035, C => n2413, D => n8025, Z => 
                           n5487);
   U1107 : AO4 port map( A => n4065, B => n8015, C => n2413, D => n8005, Z => 
                           n5488);
   U1108 : AO4 port map( A => n4066, B => n7995, C => n2413, D => n7985, Z => 
                           n5489);
   U1109 : AO4 port map( A => n4063, B => n7975, C => n2413, D => n7965, Z => 
                           n5490);
   U1110 : AO4 port map( A => n4064, B => n7955, C => n2413, D => n7945, Z => 
                           n5491);
   U1111 : AO4 port map( A => n4061, B => n7935, C => n2413, D => n7925, Z => 
                           n5492);
   U1112 : AO4 port map( A => n4062, B => n7915, C => n2413, D => n7905, Z => 
                           n5493);
   U1113 : AO4 port map( A => n4131, B => n8055, C => n2365, D => n8041, Z => 
                           n5998);
   U1114 : AO4 port map( A => n4132, B => n8035, C => n2365, D => n8021, Z => 
                           n5999);
   U1115 : AO4 port map( A => n4129, B => n8015, C => n2365, D => n8001, Z => 
                           n6000);
   U1116 : AO4 port map( A => n4130, B => n7995, C => n2365, D => n7981, Z => 
                           n6001);
   U1117 : AO4 port map( A => n4127, B => n7975, C => n2365, D => n7961, Z => 
                           n6002);
   U1118 : AO4 port map( A => n4128, B => n7955, C => n2365, D => n7941, Z => 
                           n6003);
   U1119 : AO4 port map( A => n4125, B => n7935, C => n2365, D => n7921, Z => 
                           n6004);
   U1120 : AO4 port map( A => n4126, B => n7915, C => n2365, D => n7901, Z => 
                           n6005);
   U1121 : AO4 port map( A => n4195, B => n8056, C => n2317, D => n8037, Z => 
                           n6510);
   U1122 : AO4 port map( A => n4196, B => n8036, C => n2317, D => n8017, Z => 
                           n6511);
   U1123 : AO4 port map( A => n4193, B => n8016, C => n2317, D => n7997, Z => 
                           n6512);
   U1124 : AO4 port map( A => n4194, B => n7996, C => n2317, D => n7977, Z => 
                           n6513);
   U1125 : AO4 port map( A => n4191, B => n7976, C => n2317, D => n7957, Z => 
                           n6514);
   U1126 : AO4 port map( A => n4192, B => n7956, C => n2317, D => n7937, Z => 
                           n6515);
   U1127 : AO4 port map( A => n4189, B => n7936, C => n2317, D => n7917, Z => 
                           n6516);
   U1128 : AO4 port map( A => n4190, B => n7916, C => n2317, D => n7897, Z => 
                           n6517);
   U1129 : AO4 port map( A => n4259, B => n8054, C => n6743, D => n8049, Z => 
                           n4974);
   U1131 : AO4 port map( A => n4260, B => n8034, C => n6743, D => n8029, Z => 
                           n4975);
   U1132 : AO4 port map( A => n4257, B => n8014, C => n6743, D => n8009, Z => 
                           n4976);
   U1133 : AO4 port map( A => n4258, B => n7994, C => n6743, D => n7989, Z => 
                           n4977);
   U1134 : AO4 port map( A => n4255, B => n7974, C => n6743, D => n7969, Z => 
                           n4978);
   U1135 : AO4 port map( A => n4256, B => n7954, C => n6743, D => n7949, Z => 
                           n4979);
   U1136 : AO4 port map( A => n4253, B => n7934, C => n6743, D => n7929, Z => 
                           n4980);
   U1137 : AO4 port map( A => n4254, B => n7914, C => n6743, D => n7909, Z => 
                           n4981);
   U1138 : AO4 port map( A => n4324, B => n8055, C => n2407, D => n8045, Z => 
                           n5550);
   U1139 : AO4 port map( A => n4325, B => n8035, C => n2407, D => n8025, Z => 
                           n5551);
   U1140 : AO4 port map( A => n4322, B => n8015, C => n2407, D => n8005, Z => 
                           n5552);
   U1141 : AO4 port map( A => n4323, B => n7995, C => n2407, D => n7985, Z => 
                           n5553);
   U1142 : AO4 port map( A => n4320, B => n7975, C => n2407, D => n7965, Z => 
                           n5554);
   U1143 : AO4 port map( A => n4321, B => n7955, C => n2407, D => n7945, Z => 
                           n5555);
   U1144 : AO4 port map( A => n4318, B => n7935, C => n2407, D => n7925, Z => 
                           n5556);
   U1145 : AO4 port map( A => n4319, B => n7915, C => n2407, D => n7905, Z => 
                           n5557);
   U1146 : AO4 port map( A => n4388, B => n8055, C => n2359, D => n8041, Z => 
                           n6062);
   U1147 : AO4 port map( A => n4389, B => n8035, C => n2359, D => n8021, Z => 
                           n6063);
   U1148 : AO4 port map( A => n4386, B => n8015, C => n2359, D => n8001, Z => 
                           n6064);
   U1149 : AO4 port map( A => n4387, B => n7995, C => n2359, D => n7981, Z => 
                           n6065);
   U1150 : AO4 port map( A => n4384, B => n7975, C => n2359, D => n7961, Z => 
                           n6066);
   U1151 : AO4 port map( A => n4385, B => n7955, C => n2359, D => n7941, Z => 
                           n6067);
   U1152 : AO4 port map( A => n4382, B => n7935, C => n2359, D => n7921, Z => 
                           n6068);
   U1153 : AO4 port map( A => n4383, B => n7915, C => n2359, D => n7901, Z => 
                           n6069);
   U1154 : AO4 port map( A => n4452, B => n8056, C => n2311, D => n8037, Z => 
                           n6574);
   U1155 : AO4 port map( A => n4453, B => n8036, C => n2311, D => n8017, Z => 
                           n6575);
   U1156 : AO4 port map( A => n4450, B => n8016, C => n2311, D => n7997, Z => 
                           n6576);
   U1157 : AO4 port map( A => n4451, B => n7996, C => n2311, D => n7977, Z => 
                           n6577);
   U1158 : AO4 port map( A => n4448, B => n7976, C => n2311, D => n7957, Z => 
                           n6578);
   U1159 : AO4 port map( A => n4449, B => n7956, C => n2311, D => n7937, Z => 
                           n6579);
   U1160 : AO4 port map( A => n4446, B => n7936, C => n2311, D => n7917, Z => 
                           n6580);
   U1161 : AO4 port map( A => n4447, B => n7916, C => n2311, D => n7897, Z => 
                           n6581);
   U1162 : AO4 port map( A => n4516, B => n8054, C => n6737, D => n8049, Z => 
                           n5038);
   U1163 : AO4 port map( A => n4517, B => n8034, C => n6737, D => n8029, Z => 
                           n5039);
   U1164 : AO4 port map( A => n4514, B => n8014, C => n6737, D => n8009, Z => 
                           n5040);
   U1165 : AO4 port map( A => n4515, B => n7994, C => n6737, D => n7989, Z => 
                           n5041);
   U1166 : AO4 port map( A => n4512, B => n7974, C => n6737, D => n7969, Z => 
                           n5042);
   U1167 : AO4 port map( A => n4513, B => n7954, C => n6737, D => n7949, Z => 
                           n5043);
   U1168 : AO4 port map( A => n4510, B => n7934, C => n6737, D => n7929, Z => 
                           n5044);
   U1169 : AO4 port map( A => n4511, B => n7914, C => n6737, D => n7909, Z => 
                           n5045);
   U1170 : AO2 port map( A => v_KEY32_IN_0_port, B => n266, C => 
                           v_TEMP_VECTOR_0_port, D => n271, Z => n2291);
   U1171 : AO2 port map( A => v_KEY32_IN_1_port, B => n266, C => 
                           v_TEMP_VECTOR_1_port, D => n271, Z => n2421);
   U1172 : AO2 port map( A => v_KEY32_IN_2_port, B => n266, C => 
                           v_TEMP_VECTOR_2_port, D => n271, Z => n2422);
   U1173 : AO2 port map( A => v_KEY32_IN_3_port, B => n266, C => 
                           v_TEMP_VECTOR_3_port, D => n271, Z => n2423);
   U1175 : ND4 port map( A => v_CALCULATION_CNTR_0_port, B => n8290, C => n2305
                           , D => n367, Z => n2476);
   U1176 : AO4 port map( A => n2538, B => n7894, C => n6730, D => n7888, Z => 
                           n5110);
   U1177 : AO4 port map( A => n2539, B => n7874, C => n6730, D => n7868, Z => 
                           n5111);
   U1178 : AO4 port map( A => n2536, B => n7854, C => n6730, D => n7848, Z => 
                           n5112);
   U1179 : AO4 port map( A => n2537, B => n7834, C => n6730, D => n7828, Z => 
                           n5113);
   U1180 : AO4 port map( A => n2534, B => n7814, C => n6730, D => n7808, Z => 
                           n5114);
   U1181 : AO4 port map( A => n2535, B => n7794, C => n6730, D => n7788, Z => 
                           n5115);
   U1182 : AO4 port map( A => n2532, B => n7774, C => n6730, D => n7768, Z => 
                           n5116);
   U1183 : AO4 port map( A => n2533, B => n7754, C => n6730, D => n7748, Z => 
                           n5117);
   U1184 : AO4 port map( A => n2546, B => n7734, C => n6730, D => n7728, Z => 
                           n5118);
   U1185 : AO4 port map( A => n2547, B => n7714, C => n6730, D => n7708, Z => 
                           n5119);
   U1186 : AO4 port map( A => n2544, B => n7694, C => n6730, D => n7688, Z => 
                           n5120);
   U1187 : AO4 port map( A => n2545, B => n7674, C => n6730, D => n7668, Z => 
                           n5121);
   U1188 : AO4 port map( A => n2542, B => n7654, C => n6730, D => n7648, Z => 
                           n5122);
   U1189 : AO4 port map( A => n2543, B => n7634, C => n6730, D => n7628, Z => 
                           n5123);
   U1190 : AO4 port map( A => n2540, B => n7614, C => n6729, D => n7608, Z => 
                           n5124);
   U1191 : AO4 port map( A => n2541, B => n7594, C => n6729, D => n7588, Z => 
                           n5125);
   U1192 : AO4 port map( A => n2554, B => n7574, C => n6729, D => n7568, Z => 
                           n5126);
   U1193 : AO4 port map( A => n2555, B => n7554, C => n6729, D => n7548, Z => 
                           n5127);
   U1194 : AO4 port map( A => n2552, B => n7534, C => n6729, D => n7528, Z => 
                           n5128);
   U1195 : AO4 port map( A => n2553, B => n7514, C => n6729, D => n7508, Z => 
                           n5129);
   U1196 : AO4 port map( A => n2550, B => n7494, C => n6729, D => n7488, Z => 
                           n5130);
   U1197 : AO4 port map( A => n2551, B => n7474, C => n6729, D => n7468, Z => 
                           n5131);
   U1198 : AO4 port map( A => n2548, B => n7454, C => n6729, D => n7448, Z => 
                           n5132);
   U1199 : AO4 port map( A => n2549, B => n7434, C => n6729, D => n7428, Z => 
                           n5133);
   U1200 : AO4 port map( A => n2498, B => n7414, C => n6729, D => n7408, Z => 
                           n5134);
   U1201 : AO4 port map( A => n2499, B => n7394, C => n6729, D => n7388, Z => 
                           n5135);
   U1202 : AO4 port map( A => n2496, B => n7374, C => n6729, D => n7368, Z => 
                           n5136);
   U1203 : AO4 port map( A => n2497, B => n7354, C => n6729, D => n7348, Z => 
                           n5137);
   U1204 : AO4 port map( A => n2494, B => n7334, C => n6728, D => n7328, Z => 
                           n5138);
   U1205 : AO4 port map( A => n2495, B => n7314, C => n6728, D => n7308, Z => 
                           n5139);
   U1206 : AO4 port map( A => n2492, B => n7294, C => n6728, D => n7288, Z => 
                           n5140);
   U1207 : AO4 port map( A => n2493, B => n7274, C => n6728, D => n7268, Z => 
                           n5141);
   U1208 : AO4 port map( A => n2506, B => n7254, C => n6728, D => n7248, Z => 
                           n5142);
   U1209 : AO4 port map( A => n2507, B => n7234, C => n6728, D => n7228, Z => 
                           n5143);
   U1210 : AO4 port map( A => n2504, B => n7214, C => n6728, D => n7208, Z => 
                           n5144);
   U1211 : AO4 port map( A => n2505, B => n7194, C => n6728, D => n7188, Z => 
                           n5145);
   U1212 : AO4 port map( A => n2502, B => n7174, C => n6728, D => n7168, Z => 
                           n5146);
   U1213 : AO4 port map( A => n2503, B => n7154, C => n6728, D => n7148, Z => 
                           n5147);
   U1214 : AO4 port map( A => n2500, B => n7134, C => n6728, D => n7128, Z => 
                           n5148);
   U1215 : AO4 port map( A => n2501, B => n7114, C => n6728, D => n7108, Z => 
                           n5149);
   U1216 : AO4 port map( A => n2514, B => n7094, C => n6728, D => n7088, Z => 
                           n5150);
   U1217 : AO4 port map( A => n2515, B => n7074, C => n6728, D => n7068, Z => 
                           n5151);
   U1219 : AO4 port map( A => n2512, B => n7054, C => n6727, D => n7048, Z => 
                           n5152);
   U1220 : AO4 port map( A => n2513, B => n7034, C => n6727, D => n7028, Z => 
                           n5153);
   U1221 : AO4 port map( A => n2510, B => n7014, C => n6727, D => n7008, Z => 
                           n5154);
   U1222 : AO4 port map( A => n2511, B => n6994, C => n6727, D => n6988, Z => 
                           n5155);
   U1223 : AO4 port map( A => n2508, B => n6974, C => n6727, D => n6968, Z => 
                           n5156);
   U1224 : AO4 port map( A => n2509, B => n6954, C => n6727, D => n6948, Z => 
                           n5157);
   U1225 : AO4 port map( A => n2522, B => n6934, C => n6727, D => n6928, Z => 
                           n5158);
   U1226 : AO4 port map( A => n2523, B => n6914, C => n6727, D => n6908, Z => 
                           n5159);
   U1227 : AO4 port map( A => n2520, B => n6894, C => n6727, D => n6888, Z => 
                           n5160);
   U1228 : AO4 port map( A => n2521, B => n6874, C => n6727, D => n6868, Z => 
                           n5161);
   U1229 : AO4 port map( A => n2518, B => n6854, C => n6727, D => n6848, Z => 
                           n5162);
   U1230 : AO4 port map( A => n2519, B => n6834, C => n6727, D => n6828, Z => 
                           n5163);
   U1231 : AO4 port map( A => n2516, B => n6814, C => n6727, D => n6808, Z => 
                           n5164);
   U1232 : AO4 port map( A => n2517, B => n6794, C => n6727, D => n6788, Z => 
                           n5165);
   U1233 : AO4 port map( A => n2602, B => n7895, C => n2400, D => n7884, Z => 
                           n5622);
   U1234 : AO4 port map( A => n2603, B => n7875, C => n2400, D => n7864, Z => 
                           n5623);
   U1235 : AO4 port map( A => n2600, B => n7855, C => n2400, D => n7844, Z => 
                           n5624);
   U1236 : AO4 port map( A => n2601, B => n7835, C => n2400, D => n7824, Z => 
                           n5625);
   U1237 : AO4 port map( A => n2598, B => n7815, C => n2400, D => n7804, Z => 
                           n5626);
   U1238 : AO4 port map( A => n2599, B => n7795, C => n2400, D => n7784, Z => 
                           n5627);
   U1239 : AO4 port map( A => n2596, B => n7775, C => n2400, D => n7764, Z => 
                           n5628);
   U1240 : AO4 port map( A => n2597, B => n7755, C => n2400, D => n7744, Z => 
                           n5629);
   U1241 : AO4 port map( A => n2610, B => n7735, C => n2400, D => n7724, Z => 
                           n5630);
   U1242 : AO4 port map( A => n2611, B => n7715, C => n2400, D => n7704, Z => 
                           n5631);
   U1243 : AO4 port map( A => n2608, B => n7695, C => n2400, D => n7684, Z => 
                           n5632);
   U1244 : AO4 port map( A => n2609, B => n7675, C => n2400, D => n7664, Z => 
                           n5633);
   U1245 : AO4 port map( A => n2606, B => n7655, C => n2400, D => n7644, Z => 
                           n5634);
   U1246 : AO4 port map( A => n2607, B => n7635, C => n2400, D => n7624, Z => 
                           n5635);
   U1247 : AO4 port map( A => n2604, B => n7615, C => n2399, D => n7604, Z => 
                           n5636);
   U1248 : AO4 port map( A => n2605, B => n7595, C => n2399, D => n7584, Z => 
                           n5637);
   U1249 : AO4 port map( A => n2618, B => n7575, C => n2399, D => n7564, Z => 
                           n5638);
   U1250 : AO4 port map( A => n2619, B => n7555, C => n2399, D => n7544, Z => 
                           n5639);
   U1251 : AO4 port map( A => n2616, B => n7535, C => n2399, D => n7524, Z => 
                           n5640);
   U1252 : AO4 port map( A => n2617, B => n7515, C => n2399, D => n7504, Z => 
                           n5641);
   U1253 : AO4 port map( A => n2614, B => n7495, C => n2399, D => n7484, Z => 
                           n5642);
   U1254 : AO4 port map( A => n2615, B => n7475, C => n2399, D => n7464, Z => 
                           n5643);
   U1255 : AO4 port map( A => n2612, B => n7455, C => n2399, D => n7444, Z => 
                           n5644);
   U1256 : AO4 port map( A => n2613, B => n7435, C => n2399, D => n7424, Z => 
                           n5645);
   U1257 : AO4 port map( A => n2562, B => n7415, C => n2399, D => n7404, Z => 
                           n5646);
   U1258 : AO4 port map( A => n2563, B => n7395, C => n2399, D => n7384, Z => 
                           n5647);
   U1259 : AO4 port map( A => n2560, B => n7375, C => n2399, D => n7364, Z => 
                           n5648);
   U1260 : AO4 port map( A => n2561, B => n7355, C => n2399, D => n7344, Z => 
                           n5649);
   U1261 : AO4 port map( A => n2558, B => n7335, C => n2398, D => n7324, Z => 
                           n5650);
   U1263 : AO4 port map( A => n2559, B => n7315, C => n2398, D => n7304, Z => 
                           n5651);
   U1264 : AO4 port map( A => n2556, B => n7295, C => n2398, D => n7284, Z => 
                           n5652);
   U1265 : AO4 port map( A => n2557, B => n7275, C => n2398, D => n7264, Z => 
                           n5653);
   U1266 : AO4 port map( A => n2570, B => n7255, C => n2398, D => n7244, Z => 
                           n5654);
   U1267 : AO4 port map( A => n2571, B => n7235, C => n2398, D => n7224, Z => 
                           n5655);
   U1268 : AO4 port map( A => n2568, B => n7215, C => n2398, D => n7204, Z => 
                           n5656);
   U1269 : AO4 port map( A => n2569, B => n7195, C => n2398, D => n7184, Z => 
                           n5657);
   U1270 : AO4 port map( A => n2566, B => n7175, C => n2398, D => n7164, Z => 
                           n5658);
   U1271 : AO4 port map( A => n2567, B => n7155, C => n2398, D => n7144, Z => 
                           n5659);
   U1272 : AO4 port map( A => n2564, B => n7135, C => n2398, D => n7124, Z => 
                           n5660);
   U1273 : AO4 port map( A => n2565, B => n7115, C => n2398, D => n7104, Z => 
                           n5661);
   U1274 : AO4 port map( A => n2578, B => n7095, C => n2398, D => n7084, Z => 
                           n5662);
   U1275 : AO4 port map( A => n2579, B => n7075, C => n2398, D => n7064, Z => 
                           n5663);
   U1276 : AO4 port map( A => n2576, B => n7055, C => n2397, D => n7044, Z => 
                           n5664);
   U1277 : AO4 port map( A => n2577, B => n7035, C => n2397, D => n7024, Z => 
                           n5665);
   U1278 : AO4 port map( A => n2574, B => n7015, C => n2397, D => n7004, Z => 
                           n5666);
   U1279 : AO4 port map( A => n2575, B => n6995, C => n2397, D => n6984, Z => 
                           n5667);
   U1280 : AO4 port map( A => n2572, B => n6975, C => n2397, D => n6964, Z => 
                           n5668);
   U1281 : AO4 port map( A => n2573, B => n6955, C => n2397, D => n6944, Z => 
                           n5669);
   U1282 : AO4 port map( A => n2586, B => n6935, C => n2397, D => n6924, Z => 
                           n5670);
   U1283 : AO4 port map( A => n2587, B => n6915, C => n2397, D => n6904, Z => 
                           n5671);
   U1284 : AO4 port map( A => n2584, B => n6895, C => n2397, D => n6884, Z => 
                           n5672);
   U1285 : AO4 port map( A => n2585, B => n6875, C => n2397, D => n6864, Z => 
                           n5673);
   U1286 : AO4 port map( A => n2582, B => n6855, C => n2397, D => n6844, Z => 
                           n5674);
   U1287 : AO4 port map( A => n2583, B => n6835, C => n2397, D => n6824, Z => 
                           n5675);
   U1288 : AO4 port map( A => n2580, B => n6815, C => n2397, D => n6804, Z => 
                           n5676);
   U1289 : AO4 port map( A => n2581, B => n6795, C => n2397, D => n6784, Z => 
                           n5677);
   U1290 : AO4 port map( A => n2666, B => n7895, C => n2352, D => n7880, Z => 
                           n6134);
   U1291 : AO4 port map( A => n2667, B => n7875, C => n2352, D => n7860, Z => 
                           n6135);
   U1292 : AO4 port map( A => n2664, B => n7855, C => n2352, D => n7840, Z => 
                           n6136);
   U1293 : AO4 port map( A => n2665, B => n7835, C => n2352, D => n7820, Z => 
                           n6137);
   U1294 : AO4 port map( A => n2662, B => n7815, C => n2352, D => n7800, Z => 
                           n6138);
   U1295 : AO4 port map( A => n2663, B => n7795, C => n2352, D => n7780, Z => 
                           n6139);
   U1296 : AO4 port map( A => n2660, B => n7775, C => n2352, D => n7760, Z => 
                           n6140);
   U1297 : AO4 port map( A => n2661, B => n7755, C => n2352, D => n7740, Z => 
                           n6141);
   U1298 : AO4 port map( A => n2674, B => n7735, C => n2352, D => n7720, Z => 
                           n6142);
   U1299 : AO4 port map( A => n2675, B => n7715, C => n2352, D => n7700, Z => 
                           n6143);
   U1300 : AO4 port map( A => n2672, B => n7695, C => n2352, D => n7680, Z => 
                           n6144);
   U1301 : AO4 port map( A => n2673, B => n7675, C => n2352, D => n7660, Z => 
                           n6145);
   U1302 : AO4 port map( A => n2670, B => n7655, C => n2352, D => n7640, Z => 
                           n6146);
   U1303 : AO4 port map( A => n2671, B => n7635, C => n2352, D => n7620, Z => 
                           n6147);
   U1304 : AO4 port map( A => n2668, B => n7615, C => n2351, D => n7600, Z => 
                           n6148);
   U1305 : AO4 port map( A => n2669, B => n7595, C => n2351, D => n7580, Z => 
                           n6149);
   U1307 : AO4 port map( A => n2682, B => n7575, C => n2351, D => n7560, Z => 
                           n6150);
   U1308 : AO4 port map( A => n2683, B => n7555, C => n2351, D => n7540, Z => 
                           n6151);
   U1309 : AO4 port map( A => n2680, B => n7535, C => n2351, D => n7520, Z => 
                           n6152);
   U1310 : AO4 port map( A => n2681, B => n7515, C => n2351, D => n7500, Z => 
                           n6153);
   U1311 : AO4 port map( A => n2678, B => n7495, C => n2351, D => n7480, Z => 
                           n6154);
   U1312 : AO4 port map( A => n2679, B => n7475, C => n2351, D => n7460, Z => 
                           n6155);
   U1313 : AO4 port map( A => n2676, B => n7455, C => n2351, D => n7440, Z => 
                           n6156);
   U1314 : AO4 port map( A => n2677, B => n7435, C => n2351, D => n7420, Z => 
                           n6157);
   U1315 : AO4 port map( A => n2626, B => n7415, C => n2351, D => n7400, Z => 
                           n6158);
   U1316 : AO4 port map( A => n2627, B => n7395, C => n2351, D => n7380, Z => 
                           n6159);
   U1317 : AO4 port map( A => n2624, B => n7375, C => n2351, D => n7360, Z => 
                           n6160);
   U1318 : AO4 port map( A => n2625, B => n7355, C => n2351, D => n7340, Z => 
                           n6161);
   U1319 : AO4 port map( A => n2622, B => n7335, C => n2350, D => n7320, Z => 
                           n6162);
   U1320 : AO4 port map( A => n2623, B => n7315, C => n2350, D => n7300, Z => 
                           n6163);
   U1321 : AO4 port map( A => n2620, B => n7295, C => n2350, D => n7280, Z => 
                           n6164);
   U1322 : AO4 port map( A => n2621, B => n7275, C => n2350, D => n7260, Z => 
                           n6165);
   U1323 : AO4 port map( A => n2634, B => n7255, C => n2350, D => n7240, Z => 
                           n6166);
   U1324 : AO4 port map( A => n2635, B => n7235, C => n2350, D => n7220, Z => 
                           n6167);
   U1325 : AO4 port map( A => n2632, B => n7215, C => n2350, D => n7200, Z => 
                           n6168);
   U1326 : AO4 port map( A => n2633, B => n7195, C => n2350, D => n7180, Z => 
                           n6169);
   U1327 : AO4 port map( A => n2630, B => n7175, C => n2350, D => n7160, Z => 
                           n6170);
   U1328 : AO4 port map( A => n2631, B => n7155, C => n2350, D => n7140, Z => 
                           n6171);
   U1329 : AO4 port map( A => n2628, B => n7135, C => n2350, D => n7120, Z => 
                           n6172);
   U1330 : AO4 port map( A => n2629, B => n7115, C => n2350, D => n7100, Z => 
                           n6173);
   U1331 : AO4 port map( A => n2642, B => n7095, C => n2350, D => n7080, Z => 
                           n6174);
   U1332 : AO4 port map( A => n2643, B => n7075, C => n2350, D => n7060, Z => 
                           n6175);
   U1333 : AO4 port map( A => n2640, B => n7055, C => n2349, D => n7040, Z => 
                           n6176);
   U1334 : AO4 port map( A => n2641, B => n7035, C => n2349, D => n7020, Z => 
                           n6177);
   U1335 : AO4 port map( A => n2638, B => n7015, C => n2349, D => n7000, Z => 
                           n6178);
   U1336 : AO4 port map( A => n2639, B => n6995, C => n2349, D => n6980, Z => 
                           n6179);
   U1337 : AO4 port map( A => n2636, B => n6975, C => n2349, D => n6960, Z => 
                           n6180);
   U1338 : AO4 port map( A => n2637, B => n6955, C => n2349, D => n6940, Z => 
                           n6181);
   U1339 : AO4 port map( A => n2650, B => n6935, C => n2349, D => n6920, Z => 
                           n6182);
   U1340 : AO4 port map( A => n2651, B => n6915, C => n2349, D => n6900, Z => 
                           n6183);
   U1341 : AO4 port map( A => n2648, B => n6895, C => n2349, D => n6880, Z => 
                           n6184);
   U1342 : AO4 port map( A => n2649, B => n6875, C => n2349, D => n6860, Z => 
                           n6185);
   U1343 : AO4 port map( A => n2646, B => n6855, C => n2349, D => n6840, Z => 
                           n6186);
   U1344 : AO4 port map( A => n2647, B => n6835, C => n2349, D => n6820, Z => 
                           n6187);
   U1345 : AO4 port map( A => n2644, B => n6815, C => n2349, D => n6800, Z => 
                           n6188);
   U1346 : AO4 port map( A => n2645, B => n6795, C => n2349, D => n6780, Z => 
                           n6189);
   U1347 : AO4 port map( A => n2722, B => n8054, C => n8061, D => n8052, Z => 
                           n4590);
   U1348 : AO4 port map( A => n2723, B => n8034, C => n8061, D => n8032, Z => 
                           n4591);
   U1349 : AO4 port map( A => n2720, B => n8014, C => n8061, D => n8012, Z => 
                           n4592);
   U1351 : AO4 port map( A => n2721, B => n7994, C => n8061, D => n7992, Z => 
                           n4593);
   U1352 : AO4 port map( A => n2718, B => n7974, C => n8061, D => n7972, Z => 
                           n4594);
   U1353 : AO4 port map( A => n2719, B => n7954, C => n8061, D => n7952, Z => 
                           n4595);
   U1354 : AO4 port map( A => n2716, B => n7934, C => n8061, D => n7932, Z => 
                           n4596);
   U1355 : AO4 port map( A => n2717, B => n7914, C => n8061, D => n7912, Z => 
                           n4597);
   U1356 : AO4 port map( A => n2730, B => n7894, C => n8060, D => n7892, Z => 
                           n4598);
   U1357 : AO4 port map( A => n2731, B => n7874, C => n8060, D => n7872, Z => 
                           n4599);
   U1358 : AO4 port map( A => n2728, B => n7854, C => n8060, D => n7852, Z => 
                           n4600);
   U1359 : AO4 port map( A => n2729, B => n7834, C => n8060, D => n7832, Z => 
                           n4601);
   U1360 : AO4 port map( A => n2726, B => n7814, C => n8060, D => n7812, Z => 
                           n4602);
   U1361 : AO4 port map( A => n2727, B => n7794, C => n8060, D => n7792, Z => 
                           n4603);
   U1362 : AO4 port map( A => n2724, B => n7774, C => n8060, D => n7772, Z => 
                           n4604);
   U1363 : AO4 port map( A => n2725, B => n7754, C => n8060, D => n7752, Z => 
                           n4605);
   U1364 : AO4 port map( A => n2738, B => n7734, C => n8060, D => n7732, Z => 
                           n4606);
   U1365 : AO4 port map( A => n2739, B => n7714, C => n8060, D => n7712, Z => 
                           n4607);
   U1366 : AO4 port map( A => n2736, B => n7694, C => n8060, D => n7692, Z => 
                           n4608);
   U1367 : AO4 port map( A => n2737, B => n7674, C => n8060, D => n7672, Z => 
                           n4609);
   U1368 : AO4 port map( A => n2734, B => n7654, C => n8060, D => n7652, Z => 
                           n4610);
   U1369 : AO4 port map( A => n2735, B => n7634, C => n8060, D => n7632, Z => 
                           n4611);
   U1370 : AO4 port map( A => n2732, B => n7614, C => n8059, D => n7612, Z => 
                           n4612);
   U1371 : AO4 port map( A => n2733, B => n7594, C => n8059, D => n7592, Z => 
                           n4613);
   U1372 : AO4 port map( A => n2746, B => n7574, C => n8059, D => n7572, Z => 
                           n4614);
   U1373 : AO4 port map( A => n2747, B => n7554, C => n8059, D => n7552, Z => 
                           n4615);
   U1374 : AO4 port map( A => n2744, B => n7534, C => n8059, D => n7532, Z => 
                           n4616);
   U1375 : AO4 port map( A => n2745, B => n7514, C => n8059, D => n7512, Z => 
                           n4617);
   U1376 : AO4 port map( A => n2742, B => n7494, C => n8059, D => n7492, Z => 
                           n4618);
   U1377 : AO4 port map( A => n2743, B => n7474, C => n8059, D => n7472, Z => 
                           n4619);
   U1378 : AO4 port map( A => n2740, B => n7454, C => n8059, D => n7452, Z => 
                           n4620);
   U1379 : AO4 port map( A => n2741, B => n7434, C => n8059, D => n7432, Z => 
                           n4621);
   U1380 : AO4 port map( A => n2690, B => n7414, C => n8059, D => n7412, Z => 
                           n4622);
   U1381 : AO4 port map( A => n2691, B => n7394, C => n8059, D => n7392, Z => 
                           n4623);
   U1382 : AO4 port map( A => n2688, B => n7374, C => n8059, D => n7372, Z => 
                           n4624);
   U1383 : AO4 port map( A => n2689, B => n7354, C => n8059, D => n7352, Z => 
                           n4625);
   U1384 : AO4 port map( A => n2686, B => n7334, C => n8058, D => n7332, Z => 
                           n4626);
   U1385 : AO4 port map( A => n2687, B => n7314, C => n8058, D => n7312, Z => 
                           n4627);
   U1386 : AO4 port map( A => n2684, B => n7294, C => n8058, D => n7292, Z => 
                           n4628);
   U1387 : AO4 port map( A => n2685, B => n7274, C => n8058, D => n7272, Z => 
                           n4629);
   U1388 : AO4 port map( A => n2698, B => n7254, C => n8058, D => n7252, Z => 
                           n4630);
   U1389 : AO4 port map( A => n2699, B => n7234, C => n8058, D => n7232, Z => 
                           n4631);
   U1390 : AO4 port map( A => n2696, B => n7214, C => n8058, D => n7212, Z => 
                           n4632);
   U1391 : AO4 port map( A => n2697, B => n7194, C => n8058, D => n7192, Z => 
                           n4633);
   U1392 : AO4 port map( A => n2694, B => n7174, C => n8058, D => n7172, Z => 
                           n4634);
   U1393 : AO4 port map( A => n2695, B => n7154, C => n8058, D => n7152, Z => 
                           n4635);
   U1395 : AO4 port map( A => n2692, B => n7134, C => n8058, D => n7132, Z => 
                           n4636);
   U1396 : AO4 port map( A => n2693, B => n7114, C => n8058, D => n7112, Z => 
                           n4637);
   U1397 : AO4 port map( A => n2706, B => n7094, C => n8058, D => n7092, Z => 
                           n4638);
   U1398 : AO4 port map( A => n2707, B => n7074, C => n8058, D => n7072, Z => 
                           n4639);
   U1399 : AO4 port map( A => n2704, B => n7054, C => n8057, D => n7052, Z => 
                           n4640);
   U1400 : AO4 port map( A => n2705, B => n7034, C => n8057, D => n7032, Z => 
                           n4641);
   U1401 : AO4 port map( A => n2702, B => n7014, C => n8057, D => n7012, Z => 
                           n4642);
   U1402 : AO4 port map( A => n2703, B => n6994, C => n8057, D => n6992, Z => 
                           n4643);
   U1403 : AO4 port map( A => n2700, B => n6974, C => n8057, D => n6972, Z => 
                           n4644);
   U1404 : AO4 port map( A => n2701, B => n6954, C => n8057, D => n6952, Z => 
                           n4645);
   U1405 : AO4 port map( A => n2714, B => n6934, C => n8057, D => n6932, Z => 
                           n4646);
   U1406 : AO4 port map( A => n2715, B => n6914, C => n8057, D => n6912, Z => 
                           n4647);
   U1407 : AO4 port map( A => n2712, B => n6894, C => n8057, D => n6892, Z => 
                           n4648);
   U1408 : AO4 port map( A => n2713, B => n6874, C => n8057, D => n6872, Z => 
                           n4649);
   U1409 : AO4 port map( A => n2710, B => n6854, C => n8057, D => n6852, Z => 
                           n4650);
   U1410 : AO4 port map( A => n2711, B => n6834, C => n8057, D => n6832, Z => 
                           n4651);
   U1411 : AO4 port map( A => n2708, B => n6814, C => n8057, D => n6812, Z => 
                           n4652);
   U1412 : AO4 port map( A => n2709, B => n6794, C => n8057, D => n6792, Z => 
                           n4653);
   U1413 : AO4 port map( A => n2795, B => n7894, C => n6724, D => n7888, Z => 
                           n5174);
   U1414 : AO4 port map( A => n2796, B => n7874, C => n6724, D => n7868, Z => 
                           n5175);
   U1415 : AO4 port map( A => n2793, B => n7854, C => n6724, D => n7848, Z => 
                           n5176);
   U1416 : AO4 port map( A => n2794, B => n7834, C => n6724, D => n7828, Z => 
                           n5177);
   U1417 : AO4 port map( A => n2791, B => n7814, C => n6724, D => n7808, Z => 
                           n5178);
   U1418 : AO4 port map( A => n2792, B => n7794, C => n6724, D => n7788, Z => 
                           n5179);
   U1419 : AO4 port map( A => n2789, B => n7774, C => n6724, D => n7768, Z => 
                           n5180);
   U1420 : AO4 port map( A => n2790, B => n7754, C => n6724, D => n7748, Z => 
                           n5181);
   U1421 : AO4 port map( A => n2803, B => n7734, C => n6724, D => n7728, Z => 
                           n5182);
   U1422 : AO4 port map( A => n2804, B => n7714, C => n6724, D => n7708, Z => 
                           n5183);
   U1423 : AO4 port map( A => n2801, B => n7694, C => n6724, D => n7688, Z => 
                           n5184);
   U1424 : AO4 port map( A => n2802, B => n7674, C => n6724, D => n7668, Z => 
                           n5185);
   U1425 : AO4 port map( A => n2799, B => n7654, C => n6724, D => n7648, Z => 
                           n5186);
   U1426 : AO4 port map( A => n2800, B => n7634, C => n6724, D => n7628, Z => 
                           n5187);
   U1427 : AO4 port map( A => n2797, B => n7614, C => n6723, D => n7608, Z => 
                           n5188);
   U1428 : AO4 port map( A => n2798, B => n7594, C => n6723, D => n7588, Z => 
                           n5189);
   U1429 : AO4 port map( A => n2811, B => n7574, C => n6723, D => n7568, Z => 
                           n5190);
   U1430 : AO4 port map( A => n2812, B => n7554, C => n6723, D => n7548, Z => 
                           n5191);
   U1431 : AO4 port map( A => n2809, B => n7534, C => n6723, D => n7528, Z => 
                           n5192);
   U1432 : AO4 port map( A => n2810, B => n7514, C => n6723, D => n7508, Z => 
                           n5193);
   U1433 : AO4 port map( A => n2807, B => n7494, C => n6723, D => n7488, Z => 
                           n5194);
   U1434 : AO4 port map( A => n2808, B => n7474, C => n6723, D => n7468, Z => 
                           n5195);
   U1435 : AO4 port map( A => n2805, B => n7454, C => n6723, D => n7448, Z => 
                           n5196);
   U1436 : AO4 port map( A => n2806, B => n7434, C => n6723, D => n7428, Z => 
                           n5197);
   U1437 : AO4 port map( A => n2755, B => n7414, C => n6723, D => n7408, Z => 
                           n5198);
   U1439 : AO4 port map( A => n2756, B => n7394, C => n6723, D => n7388, Z => 
                           n5199);
   U1440 : AO4 port map( A => n2753, B => n7374, C => n6723, D => n7368, Z => 
                           n5200);
   U1441 : AO4 port map( A => n2754, B => n7354, C => n6723, D => n7348, Z => 
                           n5201);
   U1442 : AO4 port map( A => n2751, B => n7334, C => n6722, D => n7328, Z => 
                           n5202);
   U1443 : AO4 port map( A => n2752, B => n7314, C => n6722, D => n7308, Z => 
                           n5203);
   U1444 : AO4 port map( A => n2749, B => n7294, C => n6722, D => n7288, Z => 
                           n5204);
   U1445 : AO4 port map( A => n2750, B => n7274, C => n6722, D => n7268, Z => 
                           n5205);
   U1446 : AO4 port map( A => n2763, B => n7254, C => n6722, D => n7248, Z => 
                           n5206);
   U1447 : AO4 port map( A => n2764, B => n7234, C => n6722, D => n7228, Z => 
                           n5207);
   U1448 : AO4 port map( A => n2761, B => n7214, C => n6722, D => n7208, Z => 
                           n5208);
   U1449 : AO4 port map( A => n2762, B => n7194, C => n6722, D => n7188, Z => 
                           n5209);
   U1450 : AO4 port map( A => n2759, B => n7174, C => n6722, D => n7168, Z => 
                           n5210);
   U1451 : AO4 port map( A => n2760, B => n7154, C => n6722, D => n7148, Z => 
                           n5211);
   U1452 : AO4 port map( A => n2757, B => n7134, C => n6722, D => n7128, Z => 
                           n5212);
   U1453 : AO4 port map( A => n2758, B => n7114, C => n6722, D => n7108, Z => 
                           n5213);
   U1454 : AO4 port map( A => n2771, B => n7094, C => n6722, D => n7088, Z => 
                           n5214);
   U1455 : AO4 port map( A => n2772, B => n7074, C => n6722, D => n7068, Z => 
                           n5215);
   U1456 : AO4 port map( A => n2769, B => n7054, C => n6721, D => n7048, Z => 
                           n5216);
   U1457 : AO4 port map( A => n2770, B => n7034, C => n6721, D => n7028, Z => 
                           n5217);
   U1458 : AO4 port map( A => n2767, B => n7014, C => n6721, D => n7008, Z => 
                           n5218);
   U1459 : AO4 port map( A => n2768, B => n6994, C => n6721, D => n6988, Z => 
                           n5219);
   U1460 : AO4 port map( A => n2765, B => n6974, C => n6721, D => n6968, Z => 
                           n5220);
   U1461 : AO4 port map( A => n2766, B => n6954, C => n6721, D => n6948, Z => 
                           n5221);
   U1462 : AO4 port map( A => n2779, B => n6934, C => n6721, D => n6928, Z => 
                           n5222);
   U1463 : AO4 port map( A => n2780, B => n6914, C => n6721, D => n6908, Z => 
                           n5223);
   U1464 : AO4 port map( A => n2777, B => n6894, C => n6721, D => n6888, Z => 
                           n5224);
   U1465 : AO4 port map( A => n2778, B => n6874, C => n6721, D => n6868, Z => 
                           n5225);
   U1466 : AO4 port map( A => n2775, B => n6854, C => n6721, D => n6848, Z => 
                           n5226);
   U1467 : AO4 port map( A => n2776, B => n6834, C => n6721, D => n6828, Z => 
                           n5227);
   U1468 : AO4 port map( A => n2773, B => n6814, C => n6721, D => n6808, Z => 
                           n5228);
   U1469 : AO4 port map( A => n2774, B => n6794, C => n6721, D => n6788, Z => 
                           n5229);
   U1470 : AO4 port map( A => n2859, B => n7895, C => n2394, D => n7884, Z => 
                           n5686);
   U1471 : AO4 port map( A => n2860, B => n7875, C => n2394, D => n7864, Z => 
                           n5687);
   U1472 : AO4 port map( A => n2857, B => n7855, C => n2394, D => n7844, Z => 
                           n5688);
   U1473 : AO4 port map( A => n2858, B => n7835, C => n2394, D => n7824, Z => 
                           n5689);
   U1474 : AO4 port map( A => n2855, B => n7815, C => n2394, D => n7804, Z => 
                           n5690);
   U1475 : AO4 port map( A => n2856, B => n7795, C => n2394, D => n7784, Z => 
                           n5691);
   U1476 : AO4 port map( A => n2853, B => n7775, C => n2394, D => n7764, Z => 
                           n5692);
   U1477 : AO4 port map( A => n2854, B => n7755, C => n2394, D => n7744, Z => 
                           n5693);
   U1478 : AO4 port map( A => n2867, B => n7735, C => n2394, D => n7724, Z => 
                           n5694);
   U1479 : AO4 port map( A => n2868, B => n7715, C => n2394, D => n7704, Z => 
                           n5695);
   U1480 : AO4 port map( A => n2865, B => n7695, C => n2394, D => n7684, Z => 
                           n5696);
   U1481 : AO4 port map( A => n2866, B => n7675, C => n2394, D => n7664, Z => 
                           n5697);
   U1483 : AO4 port map( A => n2863, B => n7655, C => n2394, D => n7644, Z => 
                           n5698);
   U1484 : AO4 port map( A => n2864, B => n7635, C => n2394, D => n7624, Z => 
                           n5699);
   U1485 : AO4 port map( A => n2861, B => n7615, C => n2393, D => n7604, Z => 
                           n5700);
   U1486 : AO4 port map( A => n2862, B => n7595, C => n2393, D => n7584, Z => 
                           n5701);
   U1487 : AO4 port map( A => n2875, B => n7575, C => n2393, D => n7564, Z => 
                           n5702);
   U1488 : AO4 port map( A => n2876, B => n7555, C => n2393, D => n7544, Z => 
                           n5703);
   U1489 : AO4 port map( A => n2873, B => n7535, C => n2393, D => n7524, Z => 
                           n5704);
   U1490 : AO4 port map( A => n2874, B => n7515, C => n2393, D => n7504, Z => 
                           n5705);
   U1491 : AO4 port map( A => n2871, B => n7495, C => n2393, D => n7484, Z => 
                           n5706);
   U1492 : AO4 port map( A => n2872, B => n7475, C => n2393, D => n7464, Z => 
                           n5707);
   U1493 : AO4 port map( A => n2869, B => n7455, C => n2393, D => n7444, Z => 
                           n5708);
   U1494 : AO4 port map( A => n2870, B => n7435, C => n2393, D => n7424, Z => 
                           n5709);
   U1495 : AO4 port map( A => n2819, B => n7415, C => n2393, D => n7404, Z => 
                           n5710);
   U1496 : AO4 port map( A => n2820, B => n7395, C => n2393, D => n7384, Z => 
                           n5711);
   U1497 : AO4 port map( A => n2817, B => n7375, C => n2393, D => n7364, Z => 
                           n5712);
   U1498 : AO4 port map( A => n2818, B => n7355, C => n2393, D => n7344, Z => 
                           n5713);
   U1499 : AO4 port map( A => n2815, B => n7335, C => n2392, D => n7324, Z => 
                           n5714);
   U1500 : AO4 port map( A => n2816, B => n7315, C => n2392, D => n7304, Z => 
                           n5715);
   U1501 : AO4 port map( A => n2813, B => n7295, C => n2392, D => n7284, Z => 
                           n5716);
   U1502 : AO4 port map( A => n2814, B => n7275, C => n2392, D => n7264, Z => 
                           n5717);
   U1503 : AO4 port map( A => n2827, B => n7255, C => n2392, D => n7244, Z => 
                           n5718);
   U1504 : AO4 port map( A => n2828, B => n7235, C => n2392, D => n7224, Z => 
                           n5719);
   U1505 : AO4 port map( A => n2825, B => n7215, C => n2392, D => n7204, Z => 
                           n5720);
   U1506 : AO4 port map( A => n2826, B => n7195, C => n2392, D => n7184, Z => 
                           n5721);
   U1507 : AO4 port map( A => n2823, B => n7175, C => n2392, D => n7164, Z => 
                           n5722);
   U1508 : AO4 port map( A => n2824, B => n7155, C => n2392, D => n7144, Z => 
                           n5723);
   U1509 : AO4 port map( A => n2821, B => n7135, C => n2392, D => n7124, Z => 
                           n5724);
   U1510 : AO4 port map( A => n2822, B => n7115, C => n2392, D => n7104, Z => 
                           n5725);
   U1511 : AO4 port map( A => n2835, B => n7095, C => n2392, D => n7084, Z => 
                           n5726);
   U1512 : AO4 port map( A => n2836, B => n7075, C => n2392, D => n7064, Z => 
                           n5727);
   U1513 : AO4 port map( A => n2833, B => n7055, C => n2391, D => n7044, Z => 
                           n5728);
   U1514 : AO4 port map( A => n2834, B => n7035, C => n2391, D => n7024, Z => 
                           n5729);
   U1515 : AO4 port map( A => n2831, B => n7015, C => n2391, D => n7004, Z => 
                           n5730);
   U1516 : AO4 port map( A => n2832, B => n6995, C => n2391, D => n6984, Z => 
                           n5731);
   U1517 : AO4 port map( A => n2829, B => n6975, C => n2391, D => n6964, Z => 
                           n5732);
   U1518 : AO4 port map( A => n2830, B => n6955, C => n2391, D => n6944, Z => 
                           n5733);
   U1519 : AO4 port map( A => n2843, B => n6935, C => n2391, D => n6924, Z => 
                           n5734);
   U1520 : AO4 port map( A => n2844, B => n6915, C => n2391, D => n6904, Z => 
                           n5735);
   U1521 : AO4 port map( A => n2841, B => n6895, C => n2391, D => n6884, Z => 
                           n5736);
   U1522 : AO4 port map( A => n2842, B => n6875, C => n2391, D => n6864, Z => 
                           n5737);
   U1523 : AO4 port map( A => n2839, B => n6855, C => n2391, D => n6844, Z => 
                           n5738);
   U1524 : AO4 port map( A => n2840, B => n6835, C => n2391, D => n6824, Z => 
                           n5739);
   U1525 : AO4 port map( A => n2837, B => n6815, C => n2391, D => n6804, Z => 
                           n5740);
   U1527 : AO4 port map( A => n2838, B => n6795, C => n2391, D => n6784, Z => 
                           n5741);
   U1528 : AO4 port map( A => n2923, B => n7895, C => n2346, D => n7880, Z => 
                           n6198);
   U1529 : AO4 port map( A => n2924, B => n7875, C => n2346, D => n7860, Z => 
                           n6199);
   U1530 : AO4 port map( A => n2921, B => n7855, C => n2346, D => n7840, Z => 
                           n6200);
   U1531 : AO4 port map( A => n2922, B => n7835, C => n2346, D => n7820, Z => 
                           n6201);
   U1532 : AO4 port map( A => n2919, B => n7815, C => n2346, D => n7800, Z => 
                           n6202);
   U1533 : AO4 port map( A => n2920, B => n7795, C => n2346, D => n7780, Z => 
                           n6203);
   U1534 : AO4 port map( A => n2917, B => n7775, C => n2346, D => n7760, Z => 
                           n6204);
   U1535 : AO4 port map( A => n2918, B => n7755, C => n2346, D => n7740, Z => 
                           n6205);
   U1536 : AO4 port map( A => n2931, B => n7735, C => n2346, D => n7720, Z => 
                           n6206);
   U1537 : AO4 port map( A => n2932, B => n7715, C => n2346, D => n7700, Z => 
                           n6207);
   U1538 : AO4 port map( A => n2929, B => n7695, C => n2346, D => n7680, Z => 
                           n6208);
   U1539 : AO4 port map( A => n2930, B => n7675, C => n2346, D => n7660, Z => 
                           n6209);
   U1540 : AO4 port map( A => n2927, B => n7655, C => n2346, D => n7640, Z => 
                           n6210);
   U1541 : AO4 port map( A => n2928, B => n7635, C => n2346, D => n7620, Z => 
                           n6211);
   U1542 : AO4 port map( A => n2925, B => n7615, C => n2345, D => n7600, Z => 
                           n6212);
   U1543 : AO4 port map( A => n2926, B => n7595, C => n2345, D => n7580, Z => 
                           n6213);
   U1544 : AO4 port map( A => n2939, B => n7575, C => n2345, D => n7560, Z => 
                           n6214);
   U1545 : AO4 port map( A => n2940, B => n7555, C => n2345, D => n7540, Z => 
                           n6215);
   U1546 : AO4 port map( A => n2937, B => n7535, C => n2345, D => n7520, Z => 
                           n6216);
   U1547 : AO4 port map( A => n2938, B => n7515, C => n2345, D => n7500, Z => 
                           n6217);
   U1548 : AO4 port map( A => n2935, B => n7495, C => n2345, D => n7480, Z => 
                           n6218);
   U1549 : AO4 port map( A => n2936, B => n7475, C => n2345, D => n7460, Z => 
                           n6219);
   U1550 : AO4 port map( A => n2933, B => n7455, C => n2345, D => n7440, Z => 
                           n6220);
   U1551 : AO4 port map( A => n2934, B => n7435, C => n2345, D => n7420, Z => 
                           n6221);
   U1552 : AO4 port map( A => n2883, B => n7415, C => n2345, D => n7400, Z => 
                           n6222);
   U1553 : AO4 port map( A => n2884, B => n7395, C => n2345, D => n7380, Z => 
                           n6223);
   U1554 : AO4 port map( A => n2881, B => n7375, C => n2345, D => n7360, Z => 
                           n6224);
   U1555 : AO4 port map( A => n2882, B => n7355, C => n2345, D => n7340, Z => 
                           n6225);
   U1556 : AO4 port map( A => n2879, B => n7335, C => n2344, D => n7320, Z => 
                           n6226);
   U1557 : AO4 port map( A => n2880, B => n7315, C => n2344, D => n7300, Z => 
                           n6227);
   U1558 : AO4 port map( A => n2877, B => n7295, C => n2344, D => n7280, Z => 
                           n6228);
   U1559 : AO4 port map( A => n2878, B => n7275, C => n2344, D => n7260, Z => 
                           n6229);
   U1560 : AO4 port map( A => n2891, B => n7255, C => n2344, D => n7240, Z => 
                           n6230);
   U1561 : AO4 port map( A => n2892, B => n7235, C => n2344, D => n7220, Z => 
                           n6231);
   U1562 : AO4 port map( A => n2889, B => n7215, C => n2344, D => n7200, Z => 
                           n6232);
   U1563 : AO4 port map( A => n2890, B => n7195, C => n2344, D => n7180, Z => 
                           n6233);
   U1564 : AO4 port map( A => n2887, B => n7175, C => n2344, D => n7160, Z => 
                           n6234);
   U1565 : AO4 port map( A => n2888, B => n7155, C => n2344, D => n7140, Z => 
                           n6235);
   U1566 : AO4 port map( A => n2885, B => n7135, C => n2344, D => n7120, Z => 
                           n6236);
   U1567 : AO4 port map( A => n2886, B => n7115, C => n2344, D => n7100, Z => 
                           n6237);
   U1568 : AO4 port map( A => n2899, B => n7095, C => n2344, D => n7080, Z => 
                           n6238);
   U1569 : AO4 port map( A => n2900, B => n7075, C => n2344, D => n7060, Z => 
                           n6239);
   U1571 : AO4 port map( A => n2897, B => n7055, C => n2343, D => n7040, Z => 
                           n6240);
   U1572 : AO4 port map( A => n2898, B => n7035, C => n2343, D => n7020, Z => 
                           n6241);
   U1573 : AO4 port map( A => n2895, B => n7015, C => n2343, D => n7000, Z => 
                           n6242);
   U1574 : AO4 port map( A => n2896, B => n6995, C => n2343, D => n6980, Z => 
                           n6243);
   U1575 : AO4 port map( A => n2893, B => n6975, C => n2343, D => n6960, Z => 
                           n6244);
   U1576 : AO4 port map( A => n2894, B => n6955, C => n2343, D => n6940, Z => 
                           n6245);
   U1577 : AO4 port map( A => n2907, B => n6935, C => n2343, D => n6920, Z => 
                           n6246);
   U1578 : AO4 port map( A => n2908, B => n6915, C => n2343, D => n6900, Z => 
                           n6247);
   U1579 : AO4 port map( A => n2905, B => n6895, C => n2343, D => n6880, Z => 
                           n6248);
   U1580 : AO4 port map( A => n2906, B => n6875, C => n2343, D => n6860, Z => 
                           n6249);
   U1581 : AO4 port map( A => n2903, B => n6855, C => n2343, D => n6840, Z => 
                           n6250);
   U1582 : AO4 port map( A => n2904, B => n6835, C => n2343, D => n6820, Z => 
                           n6251);
   U1583 : AO4 port map( A => n2901, B => n6815, C => n2343, D => n6800, Z => 
                           n6252);
   U1584 : AO4 port map( A => n2902, B => n6795, C => n2343, D => n6780, Z => 
                           n6253);
   U1585 : AO4 port map( A => n2979, B => n8054, C => n6775, D => n8052, Z => 
                           n4654);
   U1586 : AO4 port map( A => n2980, B => n8034, C => n6775, D => n8032, Z => 
                           n4655);
   U1587 : AO4 port map( A => n2977, B => n8014, C => n6775, D => n8012, Z => 
                           n4656);
   U1588 : AO4 port map( A => n2978, B => n7994, C => n6775, D => n7992, Z => 
                           n4657);
   U1589 : AO4 port map( A => n2975, B => n7974, C => n6775, D => n7972, Z => 
                           n4658);
   U1590 : AO4 port map( A => n2976, B => n7954, C => n6775, D => n7952, Z => 
                           n4659);
   U1591 : AO4 port map( A => n2973, B => n7934, C => n6775, D => n7932, Z => 
                           n4660);
   U1592 : AO4 port map( A => n2974, B => n7914, C => n6775, D => n7912, Z => 
                           n4661);
   U1593 : AO4 port map( A => n2987, B => n7894, C => n6774, D => n7892, Z => 
                           n4662);
   U1594 : AO4 port map( A => n2988, B => n7874, C => n6774, D => n7872, Z => 
                           n4663);
   U1595 : AO4 port map( A => n2985, B => n7854, C => n6774, D => n7852, Z => 
                           n4664);
   U1596 : AO4 port map( A => n2986, B => n7834, C => n6774, D => n7832, Z => 
                           n4665);
   U1597 : AO4 port map( A => n2983, B => n7814, C => n6774, D => n7812, Z => 
                           n4666);
   U1598 : AO4 port map( A => n2984, B => n7794, C => n6774, D => n7792, Z => 
                           n4667);
   U1599 : AO4 port map( A => n2981, B => n7774, C => n6774, D => n7772, Z => 
                           n4668);
   U1600 : AO4 port map( A => n2982, B => n7754, C => n6774, D => n7752, Z => 
                           n4669);
   U1601 : AO4 port map( A => n2995, B => n7734, C => n6774, D => n7732, Z => 
                           n4670);
   U1602 : AO4 port map( A => n2996, B => n7714, C => n6774, D => n7712, Z => 
                           n4671);
   U1603 : AO4 port map( A => n2993, B => n7694, C => n6774, D => n7692, Z => 
                           n4672);
   U1604 : AO4 port map( A => n2994, B => n7674, C => n6774, D => n7672, Z => 
                           n4673);
   U1605 : AO4 port map( A => n2991, B => n7654, C => n6774, D => n7652, Z => 
                           n4674);
   U1606 : AO4 port map( A => n2992, B => n7634, C => n6774, D => n7632, Z => 
                           n4675);
   U1607 : AO4 port map( A => n2989, B => n7614, C => n6773, D => n7612, Z => 
                           n4676);
   U1608 : AO4 port map( A => n2990, B => n7594, C => n6773, D => n7592, Z => 
                           n4677);
   U1609 : AO4 port map( A => n3003, B => n7574, C => n6773, D => n7572, Z => 
                           n4678);
   U1610 : AO4 port map( A => n3004, B => n7554, C => n6773, D => n7552, Z => 
                           n4679);
   U1611 : AO4 port map( A => n3001, B => n7534, C => n6773, D => n7532, Z => 
                           n4680);
   U1612 : AO4 port map( A => n3002, B => n7514, C => n6773, D => n7512, Z => 
                           n4681);
   U1613 : AO4 port map( A => n2999, B => n7494, C => n6773, D => n7492, Z => 
                           n4682);
   U1615 : AO4 port map( A => n3000, B => n7474, C => n6773, D => n7472, Z => 
                           n4683);
   U1616 : AO4 port map( A => n2997, B => n7454, C => n6773, D => n7452, Z => 
                           n4684);
   U1617 : AO4 port map( A => n2998, B => n7434, C => n6773, D => n7432, Z => 
                           n4685);
   U1618 : AO4 port map( A => n2947, B => n7414, C => n6773, D => n7412, Z => 
                           n4686);
   U1619 : AO4 port map( A => n2948, B => n7394, C => n6773, D => n7392, Z => 
                           n4687);
   U1620 : AO4 port map( A => n2945, B => n7374, C => n6773, D => n7372, Z => 
                           n4688);
   U1621 : AO4 port map( A => n2946, B => n7354, C => n6773, D => n7352, Z => 
                           n4689);
   U1622 : AO4 port map( A => n2943, B => n7334, C => n6772, D => n7332, Z => 
                           n4690);
   U1623 : AO4 port map( A => n2944, B => n7314, C => n6772, D => n7312, Z => 
                           n4691);
   U1624 : AO4 port map( A => n2941, B => n7294, C => n6772, D => n7292, Z => 
                           n4692);
   U1625 : AO4 port map( A => n2942, B => n7274, C => n6772, D => n7272, Z => 
                           n4693);
   U1626 : AO4 port map( A => n2955, B => n7254, C => n6772, D => n7252, Z => 
                           n4694);
   U1627 : AO4 port map( A => n2956, B => n7234, C => n6772, D => n7232, Z => 
                           n4695);
   U1628 : AO4 port map( A => n2953, B => n7214, C => n6772, D => n7212, Z => 
                           n4696);
   U1629 : AO4 port map( A => n2954, B => n7194, C => n6772, D => n7192, Z => 
                           n4697);
   U1630 : AO4 port map( A => n2951, B => n7174, C => n6772, D => n7172, Z => 
                           n4698);
   U1631 : AO4 port map( A => n2952, B => n7154, C => n6772, D => n7152, Z => 
                           n4699);
   U1632 : AO4 port map( A => n2949, B => n7134, C => n6772, D => n7132, Z => 
                           n4700);
   U1633 : AO4 port map( A => n2950, B => n7114, C => n6772, D => n7112, Z => 
                           n4701);
   U1634 : AO4 port map( A => n2963, B => n7094, C => n6772, D => n7092, Z => 
                           n4702);
   U1635 : AO4 port map( A => n2964, B => n7074, C => n6772, D => n7072, Z => 
                           n4703);
   U1636 : AO4 port map( A => n2961, B => n7054, C => n6771, D => n7052, Z => 
                           n4704);
   U1637 : AO4 port map( A => n2962, B => n7034, C => n6771, D => n7032, Z => 
                           n4705);
   U1638 : AO4 port map( A => n2959, B => n7014, C => n6771, D => n7012, Z => 
                           n4706);
   U1639 : AO4 port map( A => n2960, B => n6994, C => n6771, D => n6992, Z => 
                           n4707);
   U1640 : AO4 port map( A => n2957, B => n6974, C => n6771, D => n6972, Z => 
                           n4708);
   U1641 : AO4 port map( A => n2958, B => n6954, C => n6771, D => n6952, Z => 
                           n4709);
   U1642 : AO4 port map( A => n2971, B => n6934, C => n6771, D => n6932, Z => 
                           n4710);
   U1643 : AO4 port map( A => n2972, B => n6914, C => n6771, D => n6912, Z => 
                           n4711);
   U1644 : AO4 port map( A => n2969, B => n6894, C => n6771, D => n6892, Z => 
                           n4712);
   U1645 : AO4 port map( A => n2970, B => n6874, C => n6771, D => n6872, Z => 
                           n4713);
   U1646 : AO4 port map( A => n2967, B => n6854, C => n6771, D => n6852, Z => 
                           n4714);
   U1647 : AO4 port map( A => n2968, B => n6834, C => n6771, D => n6832, Z => 
                           n4715);
   U1648 : AO4 port map( A => n2965, B => n6814, C => n6771, D => n6812, Z => 
                           n4716);
   U1649 : AO4 port map( A => n2966, B => n6794, C => n6771, D => n6792, Z => 
                           n4717);
   U1650 : AO4 port map( A => n3051, B => n7894, C => n6718, D => n7887, Z => 
                           n5238);
   U1651 : AO4 port map( A => n3052, B => n7874, C => n6718, D => n7867, Z => 
                           n5239);
   U1652 : AO4 port map( A => n3049, B => n7854, C => n6718, D => n7847, Z => 
                           n5240);
   U1653 : AO4 port map( A => n3050, B => n7834, C => n6718, D => n7827, Z => 
                           n5241);
   U1654 : AO4 port map( A => n3047, B => n7814, C => n6718, D => n7807, Z => 
                           n5242);
   U1655 : AO4 port map( A => n3048, B => n7794, C => n6718, D => n7787, Z => 
                           n5243);
   U1656 : AO4 port map( A => n3045, B => n7774, C => n6718, D => n7767, Z => 
                           n5244);
   U1657 : AO4 port map( A => n3046, B => n7754, C => n6718, D => n7747, Z => 
                           n5245);
   U1659 : AO4 port map( A => n3059, B => n7734, C => n6718, D => n7727, Z => 
                           n5246);
   U1660 : AO4 port map( A => n3060, B => n7714, C => n6718, D => n7707, Z => 
                           n5247);
   U1661 : AO4 port map( A => n3057, B => n7694, C => n6718, D => n7687, Z => 
                           n5248);
   U1662 : AO4 port map( A => n3058, B => n7674, C => n6718, D => n7667, Z => 
                           n5249);
   U1663 : AO4 port map( A => n3055, B => n7654, C => n6718, D => n7647, Z => 
                           n5250);
   U1664 : AO4 port map( A => n3056, B => n7634, C => n6718, D => n7627, Z => 
                           n5251);
   U1665 : AO4 port map( A => n3053, B => n7614, C => n6717, D => n7607, Z => 
                           n5252);
   U1666 : AO4 port map( A => n3054, B => n7594, C => n6717, D => n7587, Z => 
                           n5253);
   U1667 : AO4 port map( A => n3067, B => n7574, C => n6717, D => n7567, Z => 
                           n5254);
   U1668 : AO4 port map( A => n3068, B => n7554, C => n6717, D => n7547, Z => 
                           n5255);
   U1669 : AO4 port map( A => n3065, B => n7534, C => n6717, D => n7527, Z => 
                           n5256);
   U1670 : AO4 port map( A => n3066, B => n7514, C => n6717, D => n7507, Z => 
                           n5257);
   U1671 : AO4 port map( A => n3063, B => n7494, C => n6717, D => n7487, Z => 
                           n5258);
   U1672 : AO4 port map( A => n3064, B => n7474, C => n6717, D => n7467, Z => 
                           n5259);
   U1673 : AO4 port map( A => n3061, B => n7454, C => n6717, D => n7447, Z => 
                           n5260);
   U1674 : AO4 port map( A => n3062, B => n7434, C => n6717, D => n7427, Z => 
                           n5261);
   U1675 : AO4 port map( A => n3011, B => n7414, C => n6717, D => n7407, Z => 
                           n5262);
   U1676 : AO4 port map( A => n3012, B => n7394, C => n6717, D => n7387, Z => 
                           n5263);
   U1677 : AO4 port map( A => n3009, B => n7374, C => n6717, D => n7367, Z => 
                           n5264);
   U1678 : AO4 port map( A => n3010, B => n7354, C => n6717, D => n7347, Z => 
                           n5265);
   U1679 : AO4 port map( A => n3007, B => n7334, C => n6716, D => n7327, Z => 
                           n5266);
   U1680 : AO4 port map( A => n3008, B => n7314, C => n6716, D => n7307, Z => 
                           n5267);
   U1681 : AO4 port map( A => n3005, B => n7294, C => n6716, D => n7287, Z => 
                           n5268);
   U1682 : AO4 port map( A => n3006, B => n7274, C => n6716, D => n7267, Z => 
                           n5269);
   U1683 : AO4 port map( A => n3019, B => n7254, C => n6716, D => n7247, Z => 
                           n5270);
   U1684 : AO4 port map( A => n3020, B => n7234, C => n6716, D => n7227, Z => 
                           n5271);
   U1685 : AO4 port map( A => n3017, B => n7214, C => n6716, D => n7207, Z => 
                           n5272);
   U1686 : AO4 port map( A => n3018, B => n7194, C => n6716, D => n7187, Z => 
                           n5273);
   U1687 : AO4 port map( A => n3015, B => n7174, C => n6716, D => n7167, Z => 
                           n5274);
   U1688 : AO4 port map( A => n3016, B => n7154, C => n6716, D => n7147, Z => 
                           n5275);
   U1689 : AO4 port map( A => n3013, B => n7134, C => n6716, D => n7127, Z => 
                           n5276);
   U1690 : AO4 port map( A => n3014, B => n7114, C => n6716, D => n7107, Z => 
                           n5277);
   U1691 : AO4 port map( A => n3027, B => n7094, C => n6716, D => n7087, Z => 
                           n5278);
   U1692 : AO4 port map( A => n3028, B => n7074, C => n6716, D => n7067, Z => 
                           n5279);
   U1693 : AO4 port map( A => n3025, B => n7054, C => n6658, D => n7047, Z => 
                           n5280);
   U1694 : AO4 port map( A => n3026, B => n7034, C => n6658, D => n7027, Z => 
                           n5281);
   U1695 : AO4 port map( A => n3023, B => n7014, C => n6658, D => n7007, Z => 
                           n5282);
   U1696 : AO4 port map( A => n3024, B => n6994, C => n6658, D => n6987, Z => 
                           n5283);
   U1697 : AO4 port map( A => n3021, B => n6974, C => n6658, D => n6967, Z => 
                           n5284);
   U1698 : AO4 port map( A => n3022, B => n6954, C => n6658, D => n6947, Z => 
                           n5285);
   U1699 : AO4 port map( A => n3035, B => n6934, C => n6658, D => n6927, Z => 
                           n5286);
   U1700 : AO4 port map( A => n3036, B => n6914, C => n6658, D => n6907, Z => 
                           n5287);
   U1701 : AO4 port map( A => n3033, B => n6894, C => n6658, D => n6887, Z => 
                           n5288);
   U1703 : AO4 port map( A => n3034, B => n6874, C => n6658, D => n6867, Z => 
                           n5289);
   U1704 : AO4 port map( A => n3031, B => n6854, C => n6658, D => n6847, Z => 
                           n5290);
   U1705 : AO4 port map( A => n3032, B => n6834, C => n6658, D => n6827, Z => 
                           n5291);
   U1706 : AO4 port map( A => n3029, B => n6814, C => n6658, D => n6807, Z => 
                           n5292);
   U1707 : AO4 port map( A => n3030, B => n6794, C => n6658, D => n6787, Z => 
                           n5293);
   U1708 : AO4 port map( A => n3115, B => n7895, C => n2388, D => n7883, Z => 
                           n5750);
   U1709 : AO4 port map( A => n3116, B => n7875, C => n2388, D => n7863, Z => 
                           n5751);
   U1710 : AO4 port map( A => n3113, B => n7855, C => n2388, D => n7843, Z => 
                           n5752);
   U1711 : AO4 port map( A => n3114, B => n7835, C => n2388, D => n7823, Z => 
                           n5753);
   U1712 : AO4 port map( A => n3111, B => n7815, C => n2388, D => n7803, Z => 
                           n5754);
   U1713 : AO4 port map( A => n3112, B => n7795, C => n2388, D => n7783, Z => 
                           n5755);
   U1714 : AO4 port map( A => n3109, B => n7775, C => n2388, D => n7763, Z => 
                           n5756);
   U1715 : AO4 port map( A => n3110, B => n7755, C => n2388, D => n7743, Z => 
                           n5757);
   U1716 : AO4 port map( A => n3123, B => n7735, C => n2388, D => n7723, Z => 
                           n5758);
   U1717 : AO4 port map( A => n3124, B => n7715, C => n2388, D => n7703, Z => 
                           n5759);
   U1718 : AO4 port map( A => n3121, B => n7695, C => n2388, D => n7683, Z => 
                           n5760);
   U1719 : AO4 port map( A => n3122, B => n7675, C => n2388, D => n7663, Z => 
                           n5761);
   U1720 : AO4 port map( A => n3119, B => n7655, C => n2388, D => n7643, Z => 
                           n5762);
   U1721 : AO4 port map( A => n3120, B => n7635, C => n2388, D => n7623, Z => 
                           n5763);
   U1722 : AO4 port map( A => n3117, B => n7615, C => n2387, D => n7603, Z => 
                           n5764);
   U1723 : AO4 port map( A => n3118, B => n7595, C => n2387, D => n7583, Z => 
                           n5765);
   U1724 : AO4 port map( A => n3131, B => n7575, C => n2387, D => n7563, Z => 
                           n5766);
   U1725 : AO4 port map( A => n3132, B => n7555, C => n2387, D => n7543, Z => 
                           n5767);
   U1726 : AO4 port map( A => n3129, B => n7535, C => n2387, D => n7523, Z => 
                           n5768);
   U1727 : AO4 port map( A => n3130, B => n7515, C => n2387, D => n7503, Z => 
                           n5769);
   U1728 : AO4 port map( A => n3127, B => n7495, C => n2387, D => n7483, Z => 
                           n5770);
   U1729 : AO4 port map( A => n3128, B => n7475, C => n2387, D => n7463, Z => 
                           n5771);
   U1730 : AO4 port map( A => n3125, B => n7455, C => n2387, D => n7443, Z => 
                           n5772);
   U1731 : AO4 port map( A => n3126, B => n7435, C => n2387, D => n7423, Z => 
                           n5773);
   U1732 : AO4 port map( A => n3075, B => n7415, C => n2387, D => n7403, Z => 
                           n5774);
   U1733 : AO4 port map( A => n3076, B => n7395, C => n2387, D => n7383, Z => 
                           n5775);
   U1734 : AO4 port map( A => n3073, B => n7375, C => n2387, D => n7363, Z => 
                           n5776);
   U1735 : AO4 port map( A => n3074, B => n7355, C => n2387, D => n7343, Z => 
                           n5777);
   U1736 : AO4 port map( A => n3071, B => n7335, C => n2386, D => n7323, Z => 
                           n5778);
   U1737 : AO4 port map( A => n3072, B => n7315, C => n2386, D => n7303, Z => 
                           n5779);
   U1738 : AO4 port map( A => n3069, B => n7295, C => n2386, D => n7283, Z => 
                           n5780);
   U1739 : AO4 port map( A => n3070, B => n7275, C => n2386, D => n7263, Z => 
                           n5781);
   U1740 : AO4 port map( A => n3083, B => n7255, C => n2386, D => n7243, Z => 
                           n5782);
   U1741 : AO4 port map( A => n3084, B => n7235, C => n2386, D => n7223, Z => 
                           n5783);
   U1742 : AO4 port map( A => n3081, B => n7215, C => n2386, D => n7203, Z => 
                           n5784);
   U1743 : AO4 port map( A => n3082, B => n7195, C => n2386, D => n7183, Z => 
                           n5785);
   U1744 : AO4 port map( A => n3079, B => n7175, C => n2386, D => n7163, Z => 
                           n5786);
   U1745 : AO4 port map( A => n3080, B => n7155, C => n2386, D => n7143, Z => 
                           n5787);
   U1747 : AO4 port map( A => n3077, B => n7135, C => n2386, D => n7123, Z => 
                           n5788);
   U1748 : AO4 port map( A => n3078, B => n7115, C => n2386, D => n7103, Z => 
                           n5789);
   U1749 : AO4 port map( A => n3091, B => n7095, C => n2386, D => n7083, Z => 
                           n5790);
   U1750 : AO4 port map( A => n3092, B => n7075, C => n2386, D => n7063, Z => 
                           n5791);
   U1751 : AO4 port map( A => n3089, B => n7055, C => n2385, D => n7043, Z => 
                           n5792);
   U1752 : AO4 port map( A => n3090, B => n7035, C => n2385, D => n7023, Z => 
                           n5793);
   U1753 : AO4 port map( A => n3087, B => n7015, C => n2385, D => n7003, Z => 
                           n5794);
   U1754 : AO4 port map( A => n3088, B => n6995, C => n2385, D => n6983, Z => 
                           n5795);
   U1756 : AO4 port map( A => n3085, B => n6975, C => n2385, D => n6963, Z => 
                           n5796);
   U1757 : AO4 port map( A => n3086, B => n6955, C => n2385, D => n6943, Z => 
                           n5797);
   U1758 : AO4 port map( A => n3099, B => n6935, C => n2385, D => n6923, Z => 
                           n5798);
   U1759 : AO4 port map( A => n3100, B => n6915, C => n2385, D => n6903, Z => 
                           n5799);
   U1760 : AO4 port map( A => n3097, B => n6895, C => n2385, D => n6883, Z => 
                           n5800);
   U1761 : AO4 port map( A => n3098, B => n6875, C => n2385, D => n6863, Z => 
                           n5801);
   U1763 : AO4 port map( A => n3095, B => n6855, C => n2385, D => n6843, Z => 
                           n5802);
   U1764 : AO4 port map( A => n3096, B => n6835, C => n2385, D => n6823, Z => 
                           n5803);
   U1765 : AO4 port map( A => n3093, B => n6815, C => n2385, D => n6803, Z => 
                           n5804);
   U1766 : AO4 port map( A => n3094, B => n6795, C => n2385, D => n6783, Z => 
                           n5805);
   U1767 : AO4 port map( A => n3179, B => n7895, C => n2340, D => n7879, Z => 
                           n6262);
   U1768 : AO4 port map( A => n3180, B => n7875, C => n2340, D => n7859, Z => 
                           n6263);
   U1769 : AO4 port map( A => n3177, B => n7855, C => n2340, D => n7839, Z => 
                           n6264);
   U1771 : AO4 port map( A => n3178, B => n7835, C => n2340, D => n7819, Z => 
                           n6265);
   U1772 : AO4 port map( A => n3175, B => n7815, C => n2340, D => n7799, Z => 
                           n6266);
   U1773 : AO4 port map( A => n3176, B => n7795, C => n2340, D => n7779, Z => 
                           n6267);
   U1774 : AO4 port map( A => n3173, B => n7775, C => n2340, D => n7759, Z => 
                           n6268);
   U1775 : AO4 port map( A => n3174, B => n7755, C => n2340, D => n7739, Z => 
                           n6269);
   U1776 : AO4 port map( A => n3187, B => n7735, C => n2340, D => n7719, Z => 
                           n6270);
   U1779 : AO4 port map( A => n3188, B => n7715, C => n2340, D => n7699, Z => 
                           n6271);
   U1780 : AO4 port map( A => n3185, B => n7695, C => n2340, D => n7679, Z => 
                           n6272);
   U1781 : AO4 port map( A => n3186, B => n7675, C => n2340, D => n7659, Z => 
                           n6273);
   U1782 : AO4 port map( A => n3183, B => n7655, C => n2340, D => n7639, Z => 
                           n6274);
   U1783 : AO4 port map( A => n3184, B => n7635, C => n2340, D => n7619, Z => 
                           n6275);
   U1784 : AO4 port map( A => n3181, B => n7615, C => n2339, D => n7599, Z => 
                           n6276);
   U1785 : AO4 port map( A => n3182, B => n7595, C => n2339, D => n7579, Z => 
                           n6277);
   U1787 : AO4 port map( A => n3195, B => n7575, C => n2339, D => n7559, Z => 
                           n6278);
   U1788 : AO4 port map( A => n3196, B => n7555, C => n2339, D => n7539, Z => 
                           n6279);
   U1789 : AO4 port map( A => n3193, B => n7535, C => n2339, D => n7519, Z => 
                           n6280);
   U1790 : AO4 port map( A => n3194, B => n7515, C => n2339, D => n7499, Z => 
                           n6281);
   U1791 : AO4 port map( A => n3191, B => n7495, C => n2339, D => n7479, Z => 
                           n6282);
   U1792 : AO4 port map( A => n3192, B => n7475, C => n2339, D => n7459, Z => 
                           n6283);
   U1794 : AO4 port map( A => n3189, B => n7455, C => n2339, D => n7439, Z => 
                           n6284);
   U1795 : AO4 port map( A => n3190, B => n7435, C => n2339, D => n7419, Z => 
                           n6285);
   U1796 : AO4 port map( A => n3139, B => n7415, C => n2339, D => n7399, Z => 
                           n6286);
   U1797 : AO4 port map( A => n3140, B => n7395, C => n2339, D => n7379, Z => 
                           n6287);
   U1798 : AO4 port map( A => n3137, B => n7375, C => n2339, D => n7359, Z => 
                           n6288);
   U1799 : AO4 port map( A => n3138, B => n7355, C => n2339, D => n7339, Z => 
                           n6289);
   U1800 : AO4 port map( A => n3135, B => n7335, C => n2338, D => n7319, Z => 
                           n6290);
   U1802 : AO4 port map( A => n3136, B => n7315, C => n2338, D => n7299, Z => 
                           n6291);
   U1803 : AO4 port map( A => n3133, B => n7295, C => n2338, D => n7279, Z => 
                           n6292);
   U1804 : AO4 port map( A => n3134, B => n7275, C => n2338, D => n7259, Z => 
                           n6293);
   U1805 : AO4 port map( A => n3147, B => n7255, C => n2338, D => n7239, Z => 
                           n6294);
   U1806 : AO4 port map( A => n3148, B => n7235, C => n2338, D => n7219, Z => 
                           n6295);
   U1807 : AO4 port map( A => n3145, B => n7215, C => n2338, D => n7199, Z => 
                           n6296);
   U1810 : AO4 port map( A => n3146, B => n7195, C => n2338, D => n7179, Z => 
                           n6297);
   U1811 : AO4 port map( A => n3143, B => n7175, C => n2338, D => n7159, Z => 
                           n6298);
   U1812 : AO4 port map( A => n3144, B => n7155, C => n2338, D => n7139, Z => 
                           n6299);
   U1813 : AO4 port map( A => n3141, B => n7135, C => n2338, D => n7119, Z => 
                           n6300);
   U1814 : AO4 port map( A => n3142, B => n7115, C => n2338, D => n7099, Z => 
                           n6301);
   U1815 : AO4 port map( A => n3155, B => n7095, C => n2338, D => n7079, Z => 
                           n6302);
   U1816 : AO4 port map( A => n3156, B => n7075, C => n2338, D => n7059, Z => 
                           n6303);
   U1817 : AO4 port map( A => n3153, B => n7055, C => n2337, D => n7039, Z => 
                           n6304);
   U1818 : AO4 port map( A => n3154, B => n7035, C => n2337, D => n7019, Z => 
                           n6305);
   U1820 : AO4 port map( A => n3151, B => n7015, C => n2337, D => n6999, Z => 
                           n6306);
   U1821 : AO4 port map( A => n3152, B => n6995, C => n2337, D => n6979, Z => 
                           n6307);
   U1822 : AO4 port map( A => n3149, B => n6975, C => n2337, D => n6959, Z => 
                           n6308);
   U1823 : AO4 port map( A => n3150, B => n6955, C => n2337, D => n6939, Z => 
                           n6309);
   U1824 : AO4 port map( A => n3163, B => n6935, C => n2337, D => n6919, Z => 
                           n6310);
   U1825 : AO4 port map( A => n3164, B => n6915, C => n2337, D => n6899, Z => 
                           n6311);
   U1827 : AO4 port map( A => n3161, B => n6895, C => n2337, D => n6879, Z => 
                           n6312);
   U1828 : AO4 port map( A => n3162, B => n6875, C => n2337, D => n6859, Z => 
                           n6313);
   U1829 : AO4 port map( A => n3159, B => n6855, C => n2337, D => n6839, Z => 
                           n6314);
   U1830 : AO4 port map( A => n3160, B => n6835, C => n2337, D => n6819, Z => 
                           n6315);
   U1831 : AO4 port map( A => n3157, B => n6815, C => n2337, D => n6799, Z => 
                           n6316);
   U1832 : AO4 port map( A => n3158, B => n6795, C => n2337, D => n6779, Z => 
                           n6317);
   U1833 : AO4 port map( A => n3235, B => n8054, C => n6769, D => n8051, Z => 
                           n4718);
   U1835 : AO4 port map( A => n3236, B => n8034, C => n6769, D => n8031, Z => 
                           n4719);
   U1836 : AO4 port map( A => n3233, B => n8014, C => n6769, D => n8011, Z => 
                           n4720);
   U1837 : AO4 port map( A => n3234, B => n7994, C => n6769, D => n7991, Z => 
                           n4721);
   U1838 : AO4 port map( A => n3231, B => n7974, C => n6769, D => n7971, Z => 
                           n4722);
   U1839 : AO4 port map( A => n3232, B => n7954, C => n6769, D => n7951, Z => 
                           n4723);
   U1840 : AO4 port map( A => n3229, B => n7934, C => n6769, D => n7931, Z => 
                           n4724);
   U1843 : AO4 port map( A => n3230, B => n7914, C => n6769, D => n7911, Z => 
                           n4725);
   U1844 : AO4 port map( A => n3243, B => n7894, C => n6768, D => n7891, Z => 
                           n4726);
   U1845 : AO4 port map( A => n3244, B => n7874, C => n6768, D => n7871, Z => 
                           n4727);
   U1846 : AO4 port map( A => n3241, B => n7854, C => n6768, D => n7851, Z => 
                           n4728);
   U1847 : AO4 port map( A => n3242, B => n7834, C => n6768, D => n7831, Z => 
                           n4729);
   U1848 : AO4 port map( A => n3239, B => n7814, C => n6768, D => n7811, Z => 
                           n4730);
   U1849 : AO4 port map( A => n3240, B => n7794, C => n6768, D => n7791, Z => 
                           n4731);
   U1850 : AO4 port map( A => n3237, B => n7774, C => n6768, D => n7771, Z => 
                           n4732);
   U1853 : AO4 port map( A => n3238, B => n7754, C => n6768, D => n7751, Z => 
                           n4733);
   U1854 : AO4 port map( A => n3251, B => n7734, C => n6768, D => n7731, Z => 
                           n4734);
   U1855 : AO4 port map( A => n3252, B => n7714, C => n6768, D => n7711, Z => 
                           n4735);
   U1856 : AO4 port map( A => n3249, B => n7694, C => n6768, D => n7691, Z => 
                           n4736);
   U1857 : AO4 port map( A => n3250, B => n7674, C => n6768, D => n7671, Z => 
                           n4737);
   U1858 : AO4 port map( A => n3247, B => n7654, C => n6768, D => n7651, Z => 
                           n4738);
   U1861 : AO4 port map( A => n3248, B => n7634, C => n6768, D => n7631, Z => 
                           n4739);
   U1862 : AO4 port map( A => n3245, B => n7614, C => n6767, D => n7611, Z => 
                           n4740);
   U1863 : AO4 port map( A => n3246, B => n7594, C => n6767, D => n7591, Z => 
                           n4741);
   U1864 : AO4 port map( A => n3259, B => n7574, C => n6767, D => n7571, Z => 
                           n4742);
   U1865 : AO4 port map( A => n3260, B => n7554, C => n6767, D => n7551, Z => 
                           n4743);
   U1866 : AO4 port map( A => n3257, B => n7534, C => n6767, D => n7531, Z => 
                           n4744);
   U1867 : AO4 port map( A => n3258, B => n7514, C => n6767, D => n7511, Z => 
                           n4745);
   U1868 : AO4 port map( A => n3255, B => n7494, C => n6767, D => n7491, Z => 
                           n4746);
   U1871 : AO4 port map( A => n3256, B => n7474, C => n6767, D => n7471, Z => 
                           n4747);
   U1872 : AO4 port map( A => n3253, B => n7454, C => n6767, D => n7451, Z => 
                           n4748);
   U1873 : AO4 port map( A => n3254, B => n7434, C => n6767, D => n7431, Z => 
                           n4749);
   U1875 : AO4 port map( A => n3203, B => n7414, C => n6767, D => n7411, Z => 
                           n4750);
   U1877 : AO4 port map( A => n3204, B => n7394, C => n6767, D => n7391, Z => 
                           n4751);
   U1878 : AO4 port map( A => n3201, B => n7374, C => n6767, D => n7371, Z => 
                           n4752);
   U1879 : AO4 port map( A => n3202, B => n7354, C => n6767, D => n7351, Z => 
                           n4753);
   U1881 : AO4 port map( A => n3199, B => n7334, C => n6766, D => n7331, Z => 
                           n4754);
   U1882 : AO4 port map( A => n3200, B => n7314, C => n6766, D => n7311, Z => 
                           n4755);
   U1884 : AO4 port map( A => n3197, B => n7294, C => n6766, D => n7291, Z => 
                           n4756);
   U1885 : AO4 port map( A => n3198, B => n7274, C => n6766, D => n7271, Z => 
                           n4757);
   U1888 : AO4 port map( A => n3211, B => n7254, C => n6766, D => n7251, Z => 
                           n4758);
   U1889 : AO4 port map( A => n3212, B => n7234, C => n6766, D => n7231, Z => 
                           n4759);
   U1891 : AO4 port map( A => n3209, B => n7214, C => n6766, D => n7211, Z => 
                           n4760);
   U1892 : AO4 port map( A => n3210, B => n7194, C => n6766, D => n7191, Z => 
                           n4761);
   U1893 : AO4 port map( A => n3207, B => n7174, C => n6766, D => n7171, Z => 
                           n4762);
   U1894 : AO4 port map( A => n3208, B => n7154, C => n6766, D => n7151, Z => 
                           n4763);
   U1895 : AO4 port map( A => n3205, B => n7134, C => n6766, D => n7131, Z => 
                           n4764);
   U1897 : AO4 port map( A => n3206, B => n7114, C => n6766, D => n7111, Z => 
                           n4765);
   U1898 : AO4 port map( A => n3219, B => n7094, C => n6766, D => n7091, Z => 
                           n4766);
   U1900 : AO4 port map( A => n3220, B => n7074, C => n6766, D => n7071, Z => 
                           n4767);
   U1901 : AO4 port map( A => n3217, B => n7054, C => n6765, D => n7051, Z => 
                           n4768);
   U1902 : AO4 port map( A => n3218, B => n7034, C => n6765, D => n7031, Z => 
                           n4769);
   U1904 : AO4 port map( A => n3215, B => n7014, C => n6765, D => n7011, Z => 
                           n4770);
   U1906 : AO4 port map( A => n3216, B => n6994, C => n6765, D => n6991, Z => 
                           n4771);
   U1907 : AO4 port map( A => n3213, B => n6974, C => n6765, D => n6971, Z => 
                           n4772);
   U1909 : AO4 port map( A => n3214, B => n6954, C => n6765, D => n6951, Z => 
                           n4773);
   U1910 : AO4 port map( A => n3227, B => n6934, C => n6765, D => n6931, Z => 
                           n4774);
   U1911 : AO4 port map( A => n3228, B => n6914, C => n6765, D => n6911, Z => 
                           n4775);
   U1912 : AO4 port map( A => n3225, B => n6894, C => n6765, D => n6891, Z => 
                           n4776);
   U1913 : AO4 port map( A => n3226, B => n6874, C => n6765, D => n6871, Z => 
                           n4777);
   U1914 : AO4 port map( A => n3223, B => n6854, C => n6765, D => n6851, Z => 
                           n4778);
   U1915 : AO4 port map( A => n3224, B => n6834, C => n6765, D => n6831, Z => 
                           n4779);
   U1917 : AO4 port map( A => n3221, B => n6814, C => n6765, D => n6811, Z => 
                           n4780);
   U1919 : AO4 port map( A => n3222, B => n6794, C => n6765, D => n6791, Z => 
                           n4781);
   U1920 : AO4 port map( A => n3307, B => n7894, C => n6650, D => n7887, Z => 
                           n5302);
   U1921 : AO4 port map( A => n3308, B => n7874, C => n6650, D => n7867, Z => 
                           n5303);
   U1922 : AO4 port map( A => n3305, B => n7854, C => n6650, D => n7847, Z => 
                           n5304);
   U1924 : AO4 port map( A => n3306, B => n7834, C => n6650, D => n7827, Z => 
                           n5305);
   U1925 : AO4 port map( A => n3303, B => n7814, C => n6650, D => n7807, Z => 
                           n5306);
   U1928 : AO4 port map( A => n3304, B => n7794, C => n6650, D => n7787, Z => 
                           n5307);
   U1929 : AO4 port map( A => n3301, B => n7774, C => n6650, D => n7767, Z => 
                           n5308);
   U1930 : AO4 port map( A => n3302, B => n7754, C => n6650, D => n7747, Z => 
                           n5309);
   U1931 : AO4 port map( A => n3315, B => n7734, C => n6650, D => n7727, Z => 
                           n5310);
   U1933 : AO4 port map( A => n3316, B => n7714, C => n6650, D => n7707, Z => 
                           n5311);
   U1935 : AO4 port map( A => n3313, B => n7694, C => n6650, D => n7687, Z => 
                           n5312);
   U1937 : AO4 port map( A => n3314, B => n7674, C => n6650, D => n7667, Z => 
                           n5313);
   U1939 : AO4 port map( A => n3311, B => n7654, C => n6650, D => n7647, Z => 
                           n5314);
   U1942 : AO4 port map( A => n3312, B => n7634, C => n6650, D => n7627, Z => 
                           n5315);
   U1944 : AO4 port map( A => n3309, B => n7614, C => n4543, D => n7607, Z => 
                           n5316);
   U1946 : AO4 port map( A => n3310, B => n7594, C => n4543, D => n7587, Z => 
                           n5317);
   U1947 : AO4 port map( A => n3323, B => n7574, C => n4543, D => n7567, Z => 
                           n5318);
   U1948 : AO4 port map( A => n3324, B => n7554, C => n4543, D => n7547, Z => 
                           n5319);
   U1949 : AO4 port map( A => n3321, B => n7534, C => n4543, D => n7527, Z => 
                           n5320);
   U1950 : AO4 port map( A => n3322, B => n7514, C => n4543, D => n7507, Z => 
                           n5321);
   U1952 : AO4 port map( A => n3319, B => n7494, C => n4543, D => n7487, Z => 
                           n5322);
   U1953 : AO4 port map( A => n3320, B => n7474, C => n4543, D => n7467, Z => 
                           n5323);
   U1954 : AO4 port map( A => n3317, B => n7454, C => n4543, D => n7447, Z => 
                           n5324);
   U1956 : AO4 port map( A => n3318, B => n7434, C => n4543, D => n7427, Z => 
                           n5325);
   U1958 : AO4 port map( A => n3267, B => n7414, C => n4543, D => n7407, Z => 
                           n5326);
   U1959 : AO4 port map( A => n3268, B => n7394, C => n4543, D => n7387, Z => 
                           n5327);
   U1962 : AO4 port map( A => n3265, B => n7374, C => n4543, D => n7367, Z => 
                           n5328);
   U1963 : AO4 port map( A => n3266, B => n7354, C => n4543, D => n7347, Z => 
                           n5329);
   U1964 : AO4 port map( A => n3263, B => n7334, C => n4542, D => n7327, Z => 
                           n5330);
   U1965 : AO4 port map( A => n3264, B => n7314, C => n4542, D => n7307, Z => 
                           n5331);
   U1966 : AO4 port map( A => n3261, B => n7294, C => n4542, D => n7287, Z => 
                           n5332);
   U1967 : AO4 port map( A => n3262, B => n7274, C => n4542, D => n7267, Z => 
                           n5333);
   U1968 : AO4 port map( A => n3275, B => n7254, C => n4542, D => n7247, Z => 
                           n5334);
   U1969 : AO4 port map( A => n3276, B => n7234, C => n4542, D => n7227, Z => 
                           n5335);
   U1970 : AO4 port map( A => n3273, B => n7214, C => n4542, D => n7207, Z => 
                           n5336);
   U1971 : AO4 port map( A => n3274, B => n7194, C => n4542, D => n7187, Z => 
                           n5337);
   U1973 : AO4 port map( A => n3271, B => n7174, C => n4542, D => n7167, Z => 
                           n5338);
   U1976 : AO4 port map( A => n3272, B => n7154, C => n4542, D => n7147, Z => 
                           n5339);
   U1977 : AO4 port map( A => n3269, B => n7134, C => n4542, D => n7127, Z => 
                           n5340);
   U1978 : AO4 port map( A => n3270, B => n7114, C => n4542, D => n7107, Z => 
                           n5341);
   U1979 : AO4 port map( A => n3283, B => n7094, C => n4542, D => n7087, Z => 
                           n5342);
   U1980 : AO4 port map( A => n3284, B => n7074, C => n4542, D => n7067, Z => 
                           n5343);
   U1981 : AO4 port map( A => n3281, B => n7054, C => n2490, D => n7047, Z => 
                           n5344);
   U1982 : AO4 port map( A => n3282, B => n7034, C => n2490, D => n7027, Z => 
                           n5345);
   U1983 : AO4 port map( A => n3279, B => n7014, C => n2490, D => n7007, Z => 
                           n5346);
   U1984 : AO4 port map( A => n3280, B => n6994, C => n2490, D => n6987, Z => 
                           n5347);
   U1985 : AO4 port map( A => n3277, B => n6974, C => n2490, D => n6967, Z => 
                           n5348);
   U1986 : AO4 port map( A => n3278, B => n6954, C => n2490, D => n6947, Z => 
                           n5349);
   U1987 : AO4 port map( A => n3291, B => n6934, C => n2490, D => n6927, Z => 
                           n5350);
   U1988 : AO4 port map( A => n3292, B => n6914, C => n2490, D => n6907, Z => 
                           n5351);
   U1989 : AO4 port map( A => n3289, B => n6894, C => n2490, D => n6887, Z => 
                           n5352);
   U1990 : AO4 port map( A => n3290, B => n6874, C => n2490, D => n6867, Z => 
                           n5353);
   U1992 : AO4 port map( A => n3287, B => n6854, C => n2490, D => n6847, Z => 
                           n5354);
   U1994 : AO4 port map( A => n3288, B => n6834, C => n2490, D => n6827, Z => 
                           n5355);
   U1995 : AO4 port map( A => n3285, B => n6814, C => n2490, D => n6807, Z => 
                           n5356);
   U1996 : AO4 port map( A => n3286, B => n6794, C => n2490, D => n6787, Z => 
                           n5357);
   U1997 : AO4 port map( A => n3371, B => n7895, C => n2382, D => n7883, Z => 
                           n5814);
   U1999 : AO4 port map( A => n3372, B => n7875, C => n2382, D => n7863, Z => 
                           n5815);
   U2000 : AO4 port map( A => n3369, B => n7855, C => n2382, D => n7843, Z => 
                           n5816);
   U2001 : AO4 port map( A => n3370, B => n7835, C => n2382, D => n7823, Z => 
                           n5817);
   U2002 : AO4 port map( A => n3367, B => n7815, C => n2382, D => n7803, Z => 
                           n5818);
   U2004 : AO4 port map( A => n3368, B => n7795, C => n2382, D => n7783, Z => 
                           n5819);
   U2005 : AO4 port map( A => n3365, B => n7775, C => n2382, D => n7763, Z => 
                           n5820);
   U2006 : AO4 port map( A => n3366, B => n7755, C => n2382, D => n7743, Z => 
                           n5821);
   U2008 : AO4 port map( A => n3379, B => n7735, C => n2382, D => n7723, Z => 
                           n5822);
   U2009 : AO4 port map( A => n3380, B => n7715, C => n2382, D => n7703, Z => 
                           n5823);
   U2011 : AO4 port map( A => n3377, B => n7695, C => n2382, D => n7683, Z => 
                           n5824);
   U2012 : AO4 port map( A => n3378, B => n7675, C => n2382, D => n7663, Z => 
                           n5825);
   U2013 : AO4 port map( A => n3375, B => n7655, C => n2382, D => n7643, Z => 
                           n5826);
   U2014 : AO4 port map( A => n3376, B => n7635, C => n2382, D => n7623, Z => 
                           n5827);
   U2015 : AO4 port map( A => n3373, B => n7615, C => n2381, D => n7603, Z => 
                           n5828);
   U2016 : AO4 port map( A => n3374, B => n7595, C => n2381, D => n7583, Z => 
                           n5829);
   U2017 : AO4 port map( A => n3387, B => n7575, C => n2381, D => n7563, Z => 
                           n5830);
   U2018 : AO4 port map( A => n3388, B => n7555, C => n2381, D => n7543, Z => 
                           n5831);
   U2019 : AO4 port map( A => n3385, B => n7535, C => n2381, D => n7523, Z => 
                           n5832);
   U2020 : AO4 port map( A => n3386, B => n7515, C => n2381, D => n7503, Z => 
                           n5833);
   U2021 : AO4 port map( A => n3383, B => n7495, C => n2381, D => n7483, Z => 
                           n5834);
   U2022 : AO4 port map( A => n3384, B => n7475, C => n2381, D => n7463, Z => 
                           n5835);
   U2023 : AO4 port map( A => n3381, B => n7455, C => n2381, D => n7443, Z => 
                           n5836);
   U2024 : AO4 port map( A => n3382, B => n7435, C => n2381, D => n7423, Z => 
                           n5837);
   U2025 : AO4 port map( A => n3331, B => n7415, C => n2381, D => n7403, Z => 
                           n5838);
   U2027 : AO4 port map( A => n3332, B => n7395, C => n2381, D => n7383, Z => 
                           n5839);
   U2028 : AO4 port map( A => n3329, B => n7375, C => n2381, D => n7363, Z => 
                           n5840);
   U2030 : AO4 port map( A => n3330, B => n7355, C => n2381, D => n7343, Z => 
                           n5841);
   U2031 : AO4 port map( A => n3327, B => n7335, C => n2380, D => n7323, Z => 
                           n5842);
   U2032 : AO4 port map( A => n3328, B => n7315, C => n2380, D => n7303, Z => 
                           n5843);
   U2033 : AO4 port map( A => n3325, B => n7295, C => n2380, D => n7283, Z => 
                           n5844);
   U2035 : AO4 port map( A => n3326, B => n7275, C => n2380, D => n7263, Z => 
                           n5845);
   U2036 : AO4 port map( A => n3339, B => n7255, C => n2380, D => n7243, Z => 
                           n5846);
   U2038 : AO4 port map( A => n3340, B => n7235, C => n2380, D => n7223, Z => 
                           n5847);
   U2039 : AO4 port map( A => n3337, B => n7215, C => n2380, D => n7203, Z => 
                           n5848);
   U2041 : AO4 port map( A => n3338, B => n7195, C => n2380, D => n7183, Z => 
                           n5849);
   U2043 : AO4 port map( A => n3335, B => n7175, C => n2380, D => n7163, Z => 
                           n5850);
   U2044 : AO4 port map( A => n3336, B => n7155, C => n2380, D => n7143, Z => 
                           n5851);
   U2045 : AO4 port map( A => n3333, B => n7135, C => n2380, D => n7123, Z => 
                           n5852);
   U2047 : AO4 port map( A => n3334, B => n7115, C => n2380, D => n7103, Z => 
                           n5853);
   U2048 : AO4 port map( A => n3347, B => n7095, C => n2380, D => n7083, Z => 
                           n5854);
   U2049 : AO4 port map( A => n3348, B => n7075, C => n2380, D => n7063, Z => 
                           n5855);
   U2050 : AO4 port map( A => n3345, B => n7055, C => n2379, D => n7043, Z => 
                           n5856);
   U2051 : AO4 port map( A => n3346, B => n7035, C => n2379, D => n7023, Z => 
                           n5857);
   U2052 : AO4 port map( A => n3343, B => n7015, C => n2379, D => n7003, Z => 
                           n5858);
   U2055 : AO4 port map( A => n3344, B => n6995, C => n2379, D => n6983, Z => 
                           n5859);
   U2056 : AO4 port map( A => n3341, B => n6975, C => n2379, D => n6963, Z => 
                           n5860);
   U2057 : AO4 port map( A => n3342, B => n6955, C => n2379, D => n6943, Z => 
                           n5861);
   U2059 : AO4 port map( A => n3355, B => n6935, C => n2379, D => n6923, Z => 
                           n5862);
   U2060 : AO4 port map( A => n3356, B => n6915, C => n2379, D => n6903, Z => 
                           n5863);
   U2062 : AO4 port map( A => n3353, B => n6895, C => n2379, D => n6883, Z => 
                           n5864);
   U2064 : AO4 port map( A => n3354, B => n6875, C => n2379, D => n6863, Z => 
                           n5865);
   U2065 : AO4 port map( A => n3351, B => n6855, C => n2379, D => n6843, Z => 
                           n5866);
   U2066 : AO4 port map( A => n3352, B => n6835, C => n2379, D => n6823, Z => 
                           n5867);
   U2069 : AO4 port map( A => n3349, B => n6815, C => n2379, D => n6803, Z => 
                           n5868);
   U2070 : AO4 port map( A => n3350, B => n6795, C => n2379, D => n6783, Z => 
                           n5869);
   U2071 : AO4 port map( A => n3435, B => n7895, C => n2334, D => n7879, Z => 
                           n6326);
   U2072 : AO4 port map( A => n3436, B => n7875, C => n2334, D => n7859, Z => 
                           n6327);
   U2074 : AO4 port map( A => n3433, B => n7855, C => n2334, D => n7839, Z => 
                           n6328);
   U2075 : AO4 port map( A => n3434, B => n7835, C => n2334, D => n7819, Z => 
                           n6329);
   U2076 : AO4 port map( A => n3431, B => n7815, C => n2334, D => n7799, Z => 
                           n6330);
   U2078 : AO4 port map( A => n3432, B => n7795, C => n2334, D => n7779, Z => 
                           n6331);
   U2079 : AO4 port map( A => n3429, B => n7775, C => n2334, D => n7759, Z => 
                           n6332);
   U2080 : AO4 port map( A => n3430, B => n7755, C => n2334, D => n7739, Z => 
                           n6333);
   U2081 : AO4 port map( A => n3443, B => n7735, C => n2334, D => n7719, Z => 
                           n6334);
   U2082 : AO4 port map( A => n3444, B => n7715, C => n2334, D => n7699, Z => 
                           n6335);
   U2084 : AO4 port map( A => n3441, B => n7695, C => n2334, D => n7679, Z => 
                           n6336);
   U2087 : AO4 port map( A => n3442, B => n7675, C => n2334, D => n7659, Z => 
                           n6337);
   U2089 : AO4 port map( A => n3439, B => n7655, C => n2334, D => n7639, Z => 
                           n6338);
   U2091 : AO4 port map( A => n3440, B => n7635, C => n2334, D => n7619, Z => 
                           n6339);
   U2092 : AO4 port map( A => n3437, B => n7615, C => n2333, D => n7599, Z => 
                           n6340);
   U2093 : AO4 port map( A => n3438, B => n7595, C => n2333, D => n7579, Z => 
                           n6341);
   U2094 : AO4 port map( A => n3451, B => n7575, C => n2333, D => n7559, Z => 
                           n6342);
   U2095 : AO4 port map( A => n3452, B => n7555, C => n2333, D => n7539, Z => 
                           n6343);
   U2098 : AO4 port map( A => n3449, B => n7535, C => n2333, D => n7519, Z => 
                           n6344);
   U2099 : AO4 port map( A => n3450, B => n7515, C => n2333, D => n7499, Z => 
                           n6345);
   U2103 : AO4 port map( A => n3447, B => n7495, C => n2333, D => n7479, Z => 
                           n6346);
   U2105 : AO4 port map( A => n3448, B => n7475, C => n2333, D => n7459, Z => 
                           n6347);
   U2106 : AO4 port map( A => n3445, B => n7455, C => n2333, D => n7439, Z => 
                           n6348);
   U2108 : AO4 port map( A => n3446, B => n7435, C => n2333, D => n7419, Z => 
                           n6349);
   U2109 : AO4 port map( A => n3395, B => n7415, C => n2333, D => n7399, Z => 
                           n6350);
   U2115 : AO4 port map( A => n3396, B => n7395, C => n2333, D => n7379, Z => 
                           n6351);
   U2116 : AO4 port map( A => n3393, B => n7375, C => n2333, D => n7359, Z => 
                           n6352);
   U2117 : AO4 port map( A => n3394, B => n7355, C => n2333, D => n7339, Z => 
                           n6353);
   U2121 : AO4 port map( A => n3391, B => n7335, C => n2332, D => n7319, Z => 
                           n6354);
   U2122 : AO4 port map( A => n3392, B => n7315, C => n2332, D => n7299, Z => 
                           n6355);
   U2123 : AO4 port map( A => n3389, B => n7295, C => n2332, D => n7279, Z => 
                           n6356);
   U2124 : AO4 port map( A => n3390, B => n7275, C => n2332, D => n7259, Z => 
                           n6357);
   U2125 : AO4 port map( A => n3403, B => n7255, C => n2332, D => n7239, Z => 
                           n6358);
   U2126 : AO4 port map( A => n3404, B => n7235, C => n2332, D => n7219, Z => 
                           n6359);
   U2127 : AO4 port map( A => n3401, B => n7215, C => n2332, D => n7199, Z => 
                           n6360);
   U2128 : AO4 port map( A => n3402, B => n7195, C => n2332, D => n7179, Z => 
                           n6361);
   U2130 : AO4 port map( A => n3399, B => n7175, C => n2332, D => n7159, Z => 
                           n6362);
   U2132 : AO4 port map( A => n3400, B => n7155, C => n2332, D => n7139, Z => 
                           n6363);
   U2134 : AO4 port map( A => n3397, B => n7135, C => n2332, D => n7119, Z => 
                           n6364);
   U2136 : AO4 port map( A => n3398, B => n7115, C => n2332, D => n7099, Z => 
                           n6365);
   U2137 : AO4 port map( A => n3411, B => n7095, C => n2332, D => n7079, Z => 
                           n6366);
   U2139 : AO4 port map( A => n3412, B => n7075, C => n2332, D => n7059, Z => 
                           n6367);
   U2140 : AO4 port map( A => n3409, B => n7055, C => n2331, D => n7039, Z => 
                           n6368);
   U2141 : AO4 port map( A => n3410, B => n7035, C => n2331, D => n7019, Z => 
                           n6369);
   U2143 : AO4 port map( A => n3407, B => n7015, C => n2331, D => n6999, Z => 
                           n6370);
   U2147 : AO4 port map( A => n3408, B => n6995, C => n2331, D => n6979, Z => 
                           n6371);
   U2149 : AO4 port map( A => n3405, B => n6975, C => n2331, D => n6959, Z => 
                           n6372);
   U2151 : AO4 port map( A => n3406, B => n6955, C => n2331, D => n6939, Z => 
                           n6373);
   U2153 : AO4 port map( A => n3419, B => n6935, C => n2331, D => n6919, Z => 
                           n6374);
   U2156 : AO4 port map( A => n3420, B => n6915, C => n2331, D => n6899, Z => 
                           n6375);
   U2157 : AO4 port map( A => n3417, B => n6895, C => n2331, D => n6879, Z => 
                           n6376);
   U2158 : AO4 port map( A => n3418, B => n6875, C => n2331, D => n6859, Z => 
                           n6377);
   U2160 : AO4 port map( A => n3415, B => n6855, C => n2331, D => n6839, Z => 
                           n6378);
   U2161 : AO4 port map( A => n3416, B => n6835, C => n2331, D => n6819, Z => 
                           n6379);
   U2163 : AO4 port map( A => n3413, B => n6815, C => n2331, D => n6799, Z => 
                           n6380);
   U2164 : AO4 port map( A => n3414, B => n6795, C => n2331, D => n6779, Z => 
                           n6381);
   U2168 : AO4 port map( A => n3491, B => n8054, C => n6763, D => n8051, Z => 
                           n4782);
   U2170 : AO4 port map( A => n3492, B => n8034, C => n6763, D => n8031, Z => 
                           n4783);
   U2171 : AO4 port map( A => n3489, B => n8014, C => n6763, D => n8011, Z => 
                           n4784);
   U2172 : AO4 port map( A => n3490, B => n7994, C => n6763, D => n7991, Z => 
                           n4785);
   U2175 : AO4 port map( A => n3487, B => n7974, C => n6763, D => n7971, Z => 
                           n4786);
   U2176 : AO4 port map( A => n3488, B => n7954, C => n6763, D => n7951, Z => 
                           n4787);
   U2177 : AO4 port map( A => n3485, B => n7934, C => n6763, D => n7931, Z => 
                           n4788);
   U2178 : AO4 port map( A => n3486, B => n7914, C => n6763, D => n7911, Z => 
                           n4789);
   U2179 : AO4 port map( A => n3499, B => n7894, C => n6762, D => n7891, Z => 
                           n4790);
   U2180 : AO4 port map( A => n3500, B => n7874, C => n6762, D => n7871, Z => 
                           n4791);
   U2181 : AO4 port map( A => n3497, B => n7854, C => n6762, D => n7851, Z => 
                           n4792);
   U2183 : AO4 port map( A => n3498, B => n7834, C => n6762, D => n7831, Z => 
                           n4793);
   U2184 : AO4 port map( A => n3495, B => n7814, C => n6762, D => n7811, Z => 
                           n4794);
   U2185 : AO4 port map( A => n3496, B => n7794, C => n6762, D => n7791, Z => 
                           n4795);
   U2187 : AO4 port map( A => n3493, B => n7774, C => n6762, D => n7771, Z => 
                           n4796);
   U2189 : AO4 port map( A => n3494, B => n7754, C => n6762, D => n7751, Z => 
                           n4797);
   U2191 : AO4 port map( A => n3507, B => n7734, C => n6762, D => n7731, Z => 
                           n4798);
   U2195 : AO4 port map( A => n3508, B => n7714, C => n6762, D => n7711, Z => 
                           n4799);
   U2197 : AO4 port map( A => n3505, B => n7694, C => n6762, D => n7691, Z => 
                           n4800);
   U2198 : AO4 port map( A => n3506, B => n7674, C => n6762, D => n7671, Z => 
                           n4801);
   U2199 : AO4 port map( A => n3503, B => n7654, C => n6762, D => n7651, Z => 
                           n4802);
   U2200 : AO4 port map( A => n3504, B => n7634, C => n6762, D => n7631, Z => 
                           n4803);
   U2201 : AO4 port map( A => n3501, B => n7614, C => n6761, D => n7611, Z => 
                           n4804);
   U2204 : AO4 port map( A => n3502, B => n7594, C => n6761, D => n7591, Z => 
                           n4805);
   U2206 : AO4 port map( A => n3515, B => n7574, C => n6761, D => n7571, Z => 
                           n4806);
   U2207 : AO4 port map( A => n3516, B => n7554, C => n6761, D => n7551, Z => 
                           n4807);
   U2208 : AO4 port map( A => n3513, B => n7534, C => n6761, D => n7531, Z => 
                           n4808);
   U2212 : AO4 port map( A => n3514, B => n7514, C => n6761, D => n7511, Z => 
                           n4809);
   U2214 : AO4 port map( A => n3511, B => n7494, C => n6761, D => n7491, Z => 
                           n4810);
   U2215 : AO4 port map( A => n3512, B => n7474, C => n6761, D => n7471, Z => 
                           n4811);
   U2216 : AO4 port map( A => n3509, B => n7454, C => n6761, D => n7451, Z => 
                           n4812);
   U2217 : AO4 port map( A => n3510, B => n7434, C => n6761, D => n7431, Z => 
                           n4813);
   U2220 : AO4 port map( A => n3459, B => n7414, C => n6761, D => n7411, Z => 
                           n4814);
   U2223 : AO4 port map( A => n3460, B => n7394, C => n6761, D => n7391, Z => 
                           n4815);
   U2224 : AO4 port map( A => n3457, B => n7374, C => n6761, D => n7371, Z => 
                           n4816);
   U2227 : AO4 port map( A => n3458, B => n7354, C => n6761, D => n7351, Z => 
                           n4817);
   U2228 : AO4 port map( A => n3455, B => n7334, C => n6760, D => n7331, Z => 
                           n4818);
   U2229 : AO4 port map( A => n3456, B => n7314, C => n6760, D => n7311, Z => 
                           n4819);
   U2230 : AO4 port map( A => n3453, B => n7294, C => n6760, D => n7291, Z => 
                           n4820);
   U2232 : AO4 port map( A => n3454, B => n7274, C => n6760, D => n7271, Z => 
                           n4821);
   U2235 : AO4 port map( A => n3467, B => n7254, C => n6760, D => n7251, Z => 
                           n4822);
   U2238 : AO4 port map( A => n3468, B => n7234, C => n6760, D => n7231, Z => 
                           n4823);
   U2239 : AO4 port map( A => n3465, B => n7214, C => n6760, D => n7211, Z => 
                           n4824);
   U2241 : AO4 port map( A => n3466, B => n7194, C => n6760, D => n7191, Z => 
                           n4825);
   U2246 : AO4 port map( A => n3463, B => n7174, C => n6760, D => n7171, Z => 
                           n4826);
   U2248 : AO4 port map( A => n3464, B => n7154, C => n6760, D => n7151, Z => 
                           n4827);
   U2250 : AO4 port map( A => n3461, B => n7134, C => n6760, D => n7131, Z => 
                           n4828);
   U2251 : AO4 port map( A => n3462, B => n7114, C => n6760, D => n7111, Z => 
                           n4829);
   U2256 : AO4 port map( A => n3475, B => n7094, C => n6760, D => n7091, Z => 
                           n4830);
   U2259 : AO4 port map( A => n3476, B => n7074, C => n6760, D => n7071, Z => 
                           n4831);
   U2260 : AO4 port map( A => n3473, B => n7054, C => n6759, D => n7051, Z => 
                           n4832);
   U2263 : AO4 port map( A => n3474, B => n7034, C => n6759, D => n7031, Z => 
                           n4833);
   U2266 : AO4 port map( A => n3471, B => n7014, C => n6759, D => n7011, Z => 
                           n4834);
   U2268 : AO4 port map( A => n3472, B => n6994, C => n6759, D => n6991, Z => 
                           n4835);
   U2269 : AO4 port map( A => n3469, B => n6974, C => n6759, D => n6971, Z => 
                           n4836);
   U2271 : AO4 port map( A => n3470, B => n6954, C => n6759, D => n6951, Z => 
                           n4837);
   U2273 : AO4 port map( A => n3483, B => n6934, C => n6759, D => n6931, Z => 
                           n4838);
   U2276 : AO4 port map( A => n3484, B => n6914, C => n6759, D => n6911, Z => 
                           n4839);
   U2277 : AO4 port map( A => n3481, B => n6894, C => n6759, D => n6891, Z => 
                           n4840);
   U2278 : AO4 port map( A => n3482, B => n6874, C => n6759, D => n6871, Z => 
                           n4841);
   U2281 : AO4 port map( A => n3479, B => n6854, C => n6759, D => n6851, Z => 
                           n4842);
   U2284 : AO4 port map( A => n3480, B => n6834, C => n6759, D => n6831, Z => 
                           n4843);
   U2285 : AO4 port map( A => n3477, B => n6814, C => n6759, D => n6811, Z => 
                           n4844);
   U2287 : AO4 port map( A => n3478, B => n6794, C => n6759, D => n6791, Z => 
                           n4845);
   U2288 : AO4 port map( A => n3563, B => n7894, C => n2474, D => n7886, Z => 
                           n5366);
   U2289 : AO4 port map( A => n3564, B => n7874, C => n2474, D => n7866, Z => 
                           n5367);
   U2290 : AO4 port map( A => n3561, B => n7854, C => n2474, D => n7846, Z => 
                           n5368);
   U2291 : AO4 port map( A => n3562, B => n7834, C => n2474, D => n7826, Z => 
                           n5369);
   U2292 : AO4 port map( A => n3559, B => n7814, C => n2474, D => n7806, Z => 
                           n5370);
   U2293 : AO4 port map( A => n3560, B => n7794, C => n2474, D => n7786, Z => 
                           n5371);
   U2294 : AO4 port map( A => n3557, B => n7774, C => n2474, D => n7766, Z => 
                           n5372);
   U2295 : AO4 port map( A => n3558, B => n7754, C => n2474, D => n7746, Z => 
                           n5373);
   U2298 : AO4 port map( A => n3571, B => n7734, C => n2474, D => n7726, Z => 
                           n5374);
   U2300 : AO4 port map( A => n3572, B => n7714, C => n2474, D => n7706, Z => 
                           n5375);
   U2302 : AO4 port map( A => n3569, B => n7694, C => n2474, D => n7686, Z => 
                           n5376);
   U2303 : AO4 port map( A => n3570, B => n7674, C => n2474, D => n7666, Z => 
                           n5377);
   U2304 : AO4 port map( A => n3567, B => n7654, C => n2474, D => n7646, Z => 
                           n5378);
   U2307 : AO4 port map( A => n3568, B => n7634, C => n2474, D => n7626, Z => 
                           n5379);
   U2308 : AO4 port map( A => n3565, B => n7614, C => n2473, D => n7606, Z => 
                           n5380);
   U2309 : AO4 port map( A => n3566, B => n7594, C => n2473, D => n7586, Z => 
                           n5381);
   U2311 : AO4 port map( A => n3579, B => n7574, C => n2473, D => n7566, Z => 
                           n5382);
   U2312 : AO4 port map( A => n3580, B => n7554, C => n2473, D => n7546, Z => 
                           n5383);
   U2313 : AO4 port map( A => n3577, B => n7534, C => n2473, D => n7526, Z => 
                           n5384);
   U2314 : AO4 port map( A => n3578, B => n7514, C => n2473, D => n7506, Z => 
                           n5385);
   U2316 : AO4 port map( A => n3575, B => n7494, C => n2473, D => n7486, Z => 
                           n5386);
   U2317 : AO4 port map( A => n3576, B => n7474, C => n2473, D => n7466, Z => 
                           n5387);
   U2318 : AO4 port map( A => n3573, B => n7454, C => n2473, D => n7446, Z => 
                           n5388);
   U2319 : AO4 port map( A => n3574, B => n7434, C => n2473, D => n7426, Z => 
                           n5389);
   U2321 : AO4 port map( A => n3523, B => n7414, C => n2473, D => n7406, Z => 
                           n5390);
   U2323 : AO4 port map( A => n3524, B => n7394, C => n2473, D => n7386, Z => 
                           n5391);
   U2324 : AO4 port map( A => n3521, B => n7374, C => n2473, D => n7366, Z => 
                           n5392);
   U2326 : AO4 port map( A => n3522, B => n7354, C => n2473, D => n7346, Z => 
                           n5393);
   U2327 : AO4 port map( A => n3519, B => n7334, C => n2463, D => n7326, Z => 
                           n5394);
   U2328 : AO4 port map( A => n3520, B => n7314, C => n2463, D => n7306, Z => 
                           n5395);
   U2330 : AO4 port map( A => n3517, B => n7294, C => n2463, D => n7286, Z => 
                           n5396);
   U2331 : AO4 port map( A => n3518, B => n7274, C => n2463, D => n7266, Z => 
                           n5397);
   U2332 : AO4 port map( A => n3531, B => n7254, C => n2463, D => n7246, Z => 
                           n5398);
   U2334 : AO4 port map( A => n3532, B => n7234, C => n2463, D => n7226, Z => 
                           n5399);
   U2335 : AO4 port map( A => n3529, B => n7214, C => n2463, D => n7206, Z => 
                           n5400);
   U2337 : AO4 port map( A => n3530, B => n7194, C => n2463, D => n7186, Z => 
                           n5401);
   U2339 : AO4 port map( A => n3527, B => n7174, C => n2463, D => n7166, Z => 
                           n5402);
   U2341 : AO4 port map( A => n3528, B => n7154, C => n2463, D => n7146, Z => 
                           n5403);
   U2342 : AO4 port map( A => n3525, B => n7134, C => n2463, D => n7126, Z => 
                           n5404);
   U2344 : AO4 port map( A => n3526, B => n7114, C => n2463, D => n7106, Z => 
                           n5405);
   U2345 : AO4 port map( A => n3539, B => n7094, C => n2463, D => n7086, Z => 
                           n5406);
   U2348 : AO4 port map( A => n3540, B => n7074, C => n2463, D => n7066, Z => 
                           n5407);
   U2350 : AO4 port map( A => n3537, B => n7054, C => n2461, D => n7046, Z => 
                           n5408);
   U2351 : AO4 port map( A => n3538, B => n7034, C => n2461, D => n7026, Z => 
                           n5409);
   U2352 : AO4 port map( A => n3535, B => n7014, C => n2461, D => n7006, Z => 
                           n5410);
   U2354 : AO4 port map( A => n3536, B => n6994, C => n2461, D => n6986, Z => 
                           n5411);
   U2355 : AO4 port map( A => n3533, B => n6974, C => n2461, D => n6966, Z => 
                           n5412);
   U2356 : AO4 port map( A => n3534, B => n6954, C => n2461, D => n6946, Z => 
                           n5413);
   U2357 : AO4 port map( A => n3547, B => n6934, C => n2461, D => n6926, Z => 
                           n5414);
   U2358 : AO4 port map( A => n3548, B => n6914, C => n2461, D => n6906, Z => 
                           n5415);
   U2359 : AO4 port map( A => n3545, B => n6894, C => n2461, D => n6886, Z => 
                           n5416);
   U2360 : AO4 port map( A => n3546, B => n6874, C => n2461, D => n6866, Z => 
                           n5417);
   U2361 : AO4 port map( A => n3543, B => n6854, C => n2461, D => n6846, Z => 
                           n5418);
   U2362 : AO4 port map( A => n3544, B => n6834, C => n2461, D => n6826, Z => 
                           n5419);
   U2363 : AO4 port map( A => n3541, B => n6814, C => n2461, D => n6806, Z => 
                           n5420);
   U2364 : AO4 port map( A => n3542, B => n6794, C => n2461, D => n6786, Z => 
                           n5421);
   U2365 : AO4 port map( A => n3627, B => n7895, C => n2376, D => n7882, Z => 
                           n5878);
   U2366 : AO4 port map( A => n3628, B => n7875, C => n2376, D => n7862, Z => 
                           n5879);
   U2367 : AO4 port map( A => n3625, B => n7855, C => n2376, D => n7842, Z => 
                           n5880);
   U2368 : AO4 port map( A => n3626, B => n7835, C => n2376, D => n7822, Z => 
                           n5881);
   U2369 : AO4 port map( A => n3623, B => n7815, C => n2376, D => n7802, Z => 
                           n5882);
   U2370 : AO4 port map( A => n3624, B => n7795, C => n2376, D => n7782, Z => 
                           n5883);
   U2371 : AO4 port map( A => n3621, B => n7775, C => n2376, D => n7762, Z => 
                           n5884);
   U2372 : AO4 port map( A => n3622, B => n7755, C => n2376, D => n7742, Z => 
                           n5885);
   U2373 : AO4 port map( A => n3635, B => n7735, C => n2376, D => n7722, Z => 
                           n5886);
   U2374 : AO4 port map( A => n3636, B => n7715, C => n2376, D => n7702, Z => 
                           n5887);
   U2375 : AO4 port map( A => n3633, B => n7695, C => n2376, D => n7682, Z => 
                           n5888);
   U2376 : AO4 port map( A => n3634, B => n7675, C => n2376, D => n7662, Z => 
                           n5889);
   U2377 : AO4 port map( A => n3631, B => n7655, C => n2376, D => n7642, Z => 
                           n5890);
   U2378 : AO4 port map( A => n3632, B => n7635, C => n2376, D => n7622, Z => 
                           n5891);
   U2379 : AO4 port map( A => n3629, B => n7615, C => n2375, D => n7602, Z => 
                           n5892);
   U2380 : AO4 port map( A => n3630, B => n7595, C => n2375, D => n7582, Z => 
                           n5893);
   U2381 : AO4 port map( A => n3643, B => n7575, C => n2375, D => n7562, Z => 
                           n5894);
   U2382 : AO4 port map( A => n3644, B => n7555, C => n2375, D => n7542, Z => 
                           n5895);
   U2383 : AO4 port map( A => n3641, B => n7535, C => n2375, D => n7522, Z => 
                           n5896);
   U2384 : AO4 port map( A => n3642, B => n7515, C => n2375, D => n7502, Z => 
                           n5897);
   U2385 : AO4 port map( A => n3639, B => n7495, C => n2375, D => n7482, Z => 
                           n5898);
   U2386 : AO4 port map( A => n3640, B => n7475, C => n2375, D => n7462, Z => 
                           n5899);
   U2387 : AO4 port map( A => n3637, B => n7455, C => n2375, D => n7442, Z => 
                           n5900);
   U2388 : AO4 port map( A => n3638, B => n7435, C => n2375, D => n7422, Z => 
                           n5901);
   U2389 : AO4 port map( A => n3587, B => n7415, C => n2375, D => n7402, Z => 
                           n5902);
   U2390 : AO4 port map( A => n3588, B => n7395, C => n2375, D => n7382, Z => 
                           n5903);
   U2391 : AO4 port map( A => n3585, B => n7375, C => n2375, D => n7362, Z => 
                           n5904);
   U2392 : AO4 port map( A => n3586, B => n7355, C => n2375, D => n7342, Z => 
                           n5905);
   U2393 : AO4 port map( A => n3583, B => n7335, C => n2374, D => n7322, Z => 
                           n5906);
   U2394 : AO4 port map( A => n3584, B => n7315, C => n2374, D => n7302, Z => 
                           n5907);
   U2395 : AO4 port map( A => n3581, B => n7295, C => n2374, D => n7282, Z => 
                           n5908);
   U2396 : AO4 port map( A => n3582, B => n7275, C => n2374, D => n7262, Z => 
                           n5909);
   U2397 : AO4 port map( A => n3595, B => n7255, C => n2374, D => n7242, Z => 
                           n5910);
   U2398 : AO4 port map( A => n3596, B => n7235, C => n2374, D => n7222, Z => 
                           n5911);
   U2399 : AO4 port map( A => n3593, B => n7215, C => n2374, D => n7202, Z => 
                           n5912);
   U2400 : AO4 port map( A => n3594, B => n7195, C => n2374, D => n7182, Z => 
                           n5913);
   U2401 : AO4 port map( A => n3591, B => n7175, C => n2374, D => n7162, Z => 
                           n5914);
   U2402 : AO4 port map( A => n3592, B => n7155, C => n2374, D => n7142, Z => 
                           n5915);
   U2403 : AO4 port map( A => n3589, B => n7135, C => n2374, D => n7122, Z => 
                           n5916);
   U2404 : AO4 port map( A => n3590, B => n7115, C => n2374, D => n7102, Z => 
                           n5917);
   U2405 : AO4 port map( A => n3603, B => n7095, C => n2374, D => n7082, Z => 
                           n5918);
   U2406 : AO4 port map( A => n3604, B => n7075, C => n2374, D => n7062, Z => 
                           n5919);
   U2407 : AO4 port map( A => n3601, B => n7055, C => n2373, D => n7042, Z => 
                           n5920);
   U2408 : AO4 port map( A => n3602, B => n7035, C => n2373, D => n7022, Z => 
                           n5921);
   U2409 : AO4 port map( A => n3599, B => n7015, C => n2373, D => n7002, Z => 
                           n5922);
   U2410 : AO4 port map( A => n3600, B => n6995, C => n2373, D => n6982, Z => 
                           n5923);
   U2411 : AO4 port map( A => n3597, B => n6975, C => n2373, D => n6962, Z => 
                           n5924);
   U2412 : AO4 port map( A => n3598, B => n6955, C => n2373, D => n6942, Z => 
                           n5925);
   U2413 : AO4 port map( A => n3611, B => n6935, C => n2373, D => n6922, Z => 
                           n5926);
   U2414 : AO4 port map( A => n3612, B => n6915, C => n2373, D => n6902, Z => 
                           n5927);
   U2415 : AO4 port map( A => n3609, B => n6895, C => n2373, D => n6882, Z => 
                           n5928);
   U2416 : AO4 port map( A => n3610, B => n6875, C => n2373, D => n6862, Z => 
                           n5929);
   U2417 : AO4 port map( A => n3607, B => n6855, C => n2373, D => n6842, Z => 
                           n5930);
   U2418 : AO4 port map( A => n3608, B => n6835, C => n2373, D => n6822, Z => 
                           n5931);
   U2419 : AO4 port map( A => n3605, B => n6815, C => n2373, D => n6802, Z => 
                           n5932);
   U2420 : AO4 port map( A => n3606, B => n6795, C => n2373, D => n6782, Z => 
                           n5933);
   U2421 : AO4 port map( A => n3691, B => n7896, C => n2328, D => n7878, Z => 
                           n6390);
   U2422 : AO4 port map( A => n3692, B => n7876, C => n2328, D => n7858, Z => 
                           n6391);
   U2423 : AO4 port map( A => n3689, B => n7856, C => n2328, D => n7838, Z => 
                           n6392);
   U2424 : AO4 port map( A => n3690, B => n7836, C => n2328, D => n7818, Z => 
                           n6393);
   U2425 : AO4 port map( A => n3687, B => n7816, C => n2328, D => n7798, Z => 
                           n6394);
   U2426 : AO4 port map( A => n3688, B => n7796, C => n2328, D => n7778, Z => 
                           n6395);
   U2427 : AO4 port map( A => n3685, B => n7776, C => n2328, D => n7758, Z => 
                           n6396);
   U2428 : AO4 port map( A => n3686, B => n7756, C => n2328, D => n7738, Z => 
                           n6397);
   U2429 : AO4 port map( A => n3699, B => n7736, C => n2328, D => n7718, Z => 
                           n6398);
   U2430 : AO4 port map( A => n3700, B => n7716, C => n2328, D => n7698, Z => 
                           n6399);
   U2431 : AO4 port map( A => n3697, B => n7696, C => n2328, D => n7678, Z => 
                           n6400);
   U2432 : AO4 port map( A => n3698, B => n7676, C => n2328, D => n7658, Z => 
                           n6401);
   U2433 : AO4 port map( A => n3695, B => n7656, C => n2328, D => n7638, Z => 
                           n6402);
   U2434 : AO4 port map( A => n3696, B => n7636, C => n2328, D => n7618, Z => 
                           n6403);
   U2435 : AO4 port map( A => n3693, B => n7616, C => n2327, D => n7598, Z => 
                           n6404);
   U2436 : AO4 port map( A => n3694, B => n7596, C => n2327, D => n7578, Z => 
                           n6405);
   U2437 : AO4 port map( A => n3707, B => n7576, C => n2327, D => n7558, Z => 
                           n6406);
   U2438 : AO4 port map( A => n3708, B => n7556, C => n2327, D => n7538, Z => 
                           n6407);
   U2439 : AO4 port map( A => n3705, B => n7536, C => n2327, D => n7518, Z => 
                           n6408);
   U2440 : AO4 port map( A => n3706, B => n7516, C => n2327, D => n7498, Z => 
                           n6409);
   U2441 : AO4 port map( A => n3703, B => n7496, C => n2327, D => n7478, Z => 
                           n6410);
   U2442 : AO4 port map( A => n3704, B => n7476, C => n2327, D => n7458, Z => 
                           n6411);
   U2443 : AO4 port map( A => n3701, B => n7456, C => n2327, D => n7438, Z => 
                           n6412);
   U2444 : AO4 port map( A => n3702, B => n7436, C => n2327, D => n7418, Z => 
                           n6413);
   U2445 : AO4 port map( A => n3651, B => n7416, C => n2327, D => n7398, Z => 
                           n6414);
   U2446 : AO4 port map( A => n3652, B => n7396, C => n2327, D => n7378, Z => 
                           n6415);
   U2447 : AO4 port map( A => n3649, B => n7376, C => n2327, D => n7358, Z => 
                           n6416);
   U2448 : AO4 port map( A => n3650, B => n7356, C => n2327, D => n7338, Z => 
                           n6417);
   U2449 : AO4 port map( A => n3647, B => n7336, C => n2326, D => n7318, Z => 
                           n6418);
   U2450 : AO4 port map( A => n3648, B => n7316, C => n2326, D => n7298, Z => 
                           n6419);
   U2451 : AO4 port map( A => n3645, B => n7296, C => n2326, D => n7278, Z => 
                           n6420);
   U2452 : AO4 port map( A => n3646, B => n7276, C => n2326, D => n7258, Z => 
                           n6421);
   U2453 : AO4 port map( A => n3659, B => n7256, C => n2326, D => n7238, Z => 
                           n6422);
   U2454 : AO4 port map( A => n3660, B => n7236, C => n2326, D => n7218, Z => 
                           n6423);
   U2455 : AO4 port map( A => n3657, B => n7216, C => n2326, D => n7198, Z => 
                           n6424);
   U2456 : AO4 port map( A => n3658, B => n7196, C => n2326, D => n7178, Z => 
                           n6425);
   U2457 : AO4 port map( A => n3655, B => n7176, C => n2326, D => n7158, Z => 
                           n6426);
   U2458 : AO4 port map( A => n3656, B => n7156, C => n2326, D => n7138, Z => 
                           n6427);
   U2459 : AO4 port map( A => n3653, B => n7136, C => n2326, D => n7118, Z => 
                           n6428);
   U2460 : AO4 port map( A => n3654, B => n7116, C => n2326, D => n7098, Z => 
                           n6429);
   U2461 : AO4 port map( A => n3667, B => n7096, C => n2326, D => n7078, Z => 
                           n6430);
   U2462 : AO4 port map( A => n3668, B => n7076, C => n2326, D => n7058, Z => 
                           n6431);
   U2463 : AO4 port map( A => n3665, B => n7056, C => n2325, D => n7038, Z => 
                           n6432);
   U2464 : AO4 port map( A => n3666, B => n7036, C => n2325, D => n7018, Z => 
                           n6433);
   U2465 : AO4 port map( A => n3663, B => n7016, C => n2325, D => n6998, Z => 
                           n6434);
   U2466 : AO4 port map( A => n3664, B => n6996, C => n2325, D => n6978, Z => 
                           n6435);
   U2467 : AO4 port map( A => n3661, B => n6976, C => n2325, D => n6958, Z => 
                           n6436);
   U2468 : AO4 port map( A => n3662, B => n6956, C => n2325, D => n6938, Z => 
                           n6437);
   U2469 : AO4 port map( A => n3675, B => n6936, C => n2325, D => n6918, Z => 
                           n6438);
   U2470 : AO4 port map( A => n3676, B => n6916, C => n2325, D => n6898, Z => 
                           n6439);
   U2471 : AO4 port map( A => n3673, B => n6896, C => n2325, D => n6878, Z => 
                           n6440);
   U2472 : AO4 port map( A => n3674, B => n6876, C => n2325, D => n6858, Z => 
                           n6441);
   U2473 : AO4 port map( A => n3671, B => n6856, C => n2325, D => n6838, Z => 
                           n6442);
   U2474 : AO4 port map( A => n3672, B => n6836, C => n2325, D => n6818, Z => 
                           n6443);
   U2475 : AO4 port map( A => n3669, B => n6816, C => n2325, D => n6798, Z => 
                           n6444);
   U2476 : AO4 port map( A => n3670, B => n6796, C => n2325, D => n6778, Z => 
                           n6445);
   U2477 : AO4 port map( A => n3755, B => n7894, C => n6756, D => n7890, Z => 
                           n4854);
   U2478 : AO4 port map( A => n3756, B => n7874, C => n6756, D => n7870, Z => 
                           n4855);
   U2479 : AO4 port map( A => n3753, B => n7854, C => n6756, D => n7850, Z => 
                           n4856);
   U2480 : AO4 port map( A => n3754, B => n7834, C => n6756, D => n7830, Z => 
                           n4857);
   U2481 : AO4 port map( A => n3751, B => n7814, C => n6756, D => n7810, Z => 
                           n4858);
   U2482 : AO4 port map( A => n3752, B => n7794, C => n6756, D => n7790, Z => 
                           n4859);
   U2483 : AO4 port map( A => n3749, B => n7774, C => n6756, D => n7770, Z => 
                           n4860);
   U2484 : AO4 port map( A => n3750, B => n7754, C => n6756, D => n7750, Z => 
                           n4861);
   U2485 : AO4 port map( A => n3763, B => n7734, C => n6756, D => n7730, Z => 
                           n4862);
   U2486 : AO4 port map( A => n3764, B => n7714, C => n6756, D => n7710, Z => 
                           n4863);
   U2487 : AO4 port map( A => n3761, B => n7694, C => n6756, D => n7690, Z => 
                           n4864);
   U2488 : AO4 port map( A => n3762, B => n7674, C => n6756, D => n7670, Z => 
                           n4865);
   U2489 : AO4 port map( A => n3759, B => n7654, C => n6756, D => n7650, Z => 
                           n4866);
   U2490 : AO4 port map( A => n3760, B => n7634, C => n6756, D => n7630, Z => 
                           n4867);
   U2491 : AO4 port map( A => n3757, B => n7614, C => n6755, D => n7610, Z => 
                           n4868);
   U2492 : AO4 port map( A => n3758, B => n7594, C => n6755, D => n7590, Z => 
                           n4869);
   U2493 : AO4 port map( A => n3771, B => n7574, C => n6755, D => n7570, Z => 
                           n4870);
   U2494 : AO4 port map( A => n3772, B => n7554, C => n6755, D => n7550, Z => 
                           n4871);
   U2495 : AO4 port map( A => n3769, B => n7534, C => n6755, D => n7530, Z => 
                           n4872);
   U2496 : AO4 port map( A => n3770, B => n7514, C => n6755, D => n7510, Z => 
                           n4873);
   U2497 : AO4 port map( A => n3767, B => n7494, C => n6755, D => n7490, Z => 
                           n4874);
   U2498 : AO4 port map( A => n3768, B => n7474, C => n6755, D => n7470, Z => 
                           n4875);
   U2499 : AO4 port map( A => n3765, B => n7454, C => n6755, D => n7450, Z => 
                           n4876);
   U2500 : AO4 port map( A => n3766, B => n7434, C => n6755, D => n7430, Z => 
                           n4877);
   U2501 : AO4 port map( A => n3715, B => n7414, C => n6755, D => n7410, Z => 
                           n4878);
   U2502 : AO4 port map( A => n3716, B => n7394, C => n6755, D => n7390, Z => 
                           n4879);
   U2503 : AO4 port map( A => n3713, B => n7374, C => n6755, D => n7370, Z => 
                           n4880);
   U2504 : AO4 port map( A => n3714, B => n7354, C => n6755, D => n7350, Z => 
                           n4881);
   U2505 : AO4 port map( A => n3711, B => n7334, C => n6754, D => n7330, Z => 
                           n4882);
   U2506 : AO4 port map( A => n3712, B => n7314, C => n6754, D => n7310, Z => 
                           n4883);
   U2507 : AO4 port map( A => n3709, B => n7294, C => n6754, D => n7290, Z => 
                           n4884);
   U2508 : AO4 port map( A => n3710, B => n7274, C => n6754, D => n7270, Z => 
                           n4885);
   U2509 : AO4 port map( A => n3723, B => n7254, C => n6754, D => n7250, Z => 
                           n4886);
   U2510 : AO4 port map( A => n3724, B => n7234, C => n6754, D => n7230, Z => 
                           n4887);
   U2511 : AO4 port map( A => n3721, B => n7214, C => n6754, D => n7210, Z => 
                           n4888);
   U2512 : AO4 port map( A => n3722, B => n7194, C => n6754, D => n7190, Z => 
                           n4889);
   U2513 : AO4 port map( A => n3719, B => n7174, C => n6754, D => n7170, Z => 
                           n4890);
   U2514 : AO4 port map( A => n3720, B => n7154, C => n6754, D => n7150, Z => 
                           n4891);
   U2515 : AO4 port map( A => n3717, B => n7134, C => n6754, D => n7130, Z => 
                           n4892);
   U2516 : AO4 port map( A => n3718, B => n7114, C => n6754, D => n7110, Z => 
                           n4893);
   U2517 : AO4 port map( A => n3731, B => n7094, C => n6754, D => n7090, Z => 
                           n4894);
   U2518 : AO4 port map( A => n3732, B => n7074, C => n6754, D => n7070, Z => 
                           n4895);
   U2519 : AO4 port map( A => n3729, B => n7054, C => n6753, D => n7050, Z => 
                           n4896);
   U2520 : AO4 port map( A => n3730, B => n7034, C => n6753, D => n7030, Z => 
                           n4897);
   U2521 : AO4 port map( A => n3727, B => n7014, C => n6753, D => n7010, Z => 
                           n4898);
   U2522 : AO4 port map( A => n3728, B => n6994, C => n6753, D => n6990, Z => 
                           n4899);
   U2523 : AO4 port map( A => n3725, B => n6974, C => n6753, D => n6970, Z => 
                           n4900);
   U2524 : AO4 port map( A => n3726, B => n6954, C => n6753, D => n6950, Z => 
                           n4901);
   U2525 : AO4 port map( A => n3739, B => n6934, C => n6753, D => n6930, Z => 
                           n4902);
   U2526 : AO4 port map( A => n3740, B => n6914, C => n6753, D => n6910, Z => 
                           n4903);
   U2527 : AO4 port map( A => n3737, B => n6894, C => n6753, D => n6890, Z => 
                           n4904);
   U2528 : AO4 port map( A => n3738, B => n6874, C => n6753, D => n6870, Z => 
                           n4905);
   U2529 : AO4 port map( A => n3735, B => n6854, C => n6753, D => n6850, Z => 
                           n4906);
   U2530 : AO4 port map( A => n3736, B => n6834, C => n6753, D => n6830, Z => 
                           n4907);
   U2531 : AO4 port map( A => n3733, B => n6814, C => n6753, D => n6810, Z => 
                           n4908);
   U2532 : AO4 port map( A => n3734, B => n6794, C => n6753, D => n6790, Z => 
                           n4909);
   U2533 : AO4 port map( A => n3819, B => n7894, C => n2418, D => n7886, Z => 
                           n5430);
   U2534 : AO4 port map( A => n3820, B => n7874, C => n2418, D => n7866, Z => 
                           n5431);
   U2535 : AO4 port map( A => n3817, B => n7854, C => n2418, D => n7846, Z => 
                           n5432);
   U2536 : AO4 port map( A => n3818, B => n7834, C => n2418, D => n7826, Z => 
                           n5433);
   U2537 : AO4 port map( A => n3815, B => n7814, C => n2418, D => n7806, Z => 
                           n5434);
   U2538 : AO4 port map( A => n3816, B => n7794, C => n2418, D => n7786, Z => 
                           n5435);
   U2539 : AO4 port map( A => n3813, B => n7774, C => n2418, D => n7766, Z => 
                           n5436);
   U2540 : AO4 port map( A => n3814, B => n7754, C => n2418, D => n7746, Z => 
                           n5437);
   U2541 : AO4 port map( A => n3827, B => n7734, C => n2418, D => n7726, Z => 
                           n5438);
   U2542 : AO4 port map( A => n3828, B => n7714, C => n2418, D => n7706, Z => 
                           n5439);
   U2543 : AO4 port map( A => n3825, B => n7694, C => n2418, D => n7686, Z => 
                           n5440);
   U2544 : AO4 port map( A => n3826, B => n7674, C => n2418, D => n7666, Z => 
                           n5441);
   U2545 : AO4 port map( A => n3823, B => n7654, C => n2418, D => n7646, Z => 
                           n5442);
   U2546 : AO4 port map( A => n3824, B => n7634, C => n2418, D => n7626, Z => 
                           n5443);
   U2547 : AO4 port map( A => n3821, B => n7614, C => n2417, D => n7606, Z => 
                           n5444);
   U2548 : AO4 port map( A => n3822, B => n7594, C => n2417, D => n7586, Z => 
                           n5445);
   U2549 : AO4 port map( A => n3835, B => n7574, C => n2417, D => n7566, Z => 
                           n5446);
   U2550 : AO4 port map( A => n3836, B => n7554, C => n2417, D => n7546, Z => 
                           n5447);
   U2551 : AO4 port map( A => n3833, B => n7534, C => n2417, D => n7526, Z => 
                           n5448);
   U2552 : AO4 port map( A => n3834, B => n7514, C => n2417, D => n7506, Z => 
                           n5449);
   U2553 : AO4 port map( A => n3831, B => n7494, C => n2417, D => n7486, Z => 
                           n5450);
   U2554 : AO4 port map( A => n3832, B => n7474, C => n2417, D => n7466, Z => 
                           n5451);
   U2555 : AO4 port map( A => n3829, B => n7454, C => n2417, D => n7446, Z => 
                           n5452);
   U2556 : AO4 port map( A => n3830, B => n7434, C => n2417, D => n7426, Z => 
                           n5453);
   U2557 : AO4 port map( A => n3779, B => n7414, C => n2417, D => n7406, Z => 
                           n5454);
   U2558 : AO4 port map( A => n3780, B => n7394, C => n2417, D => n7386, Z => 
                           n5455);
   U2559 : AO4 port map( A => n3777, B => n7374, C => n2417, D => n7366, Z => 
                           n5456);
   U2560 : AO4 port map( A => n3778, B => n7354, C => n2417, D => n7346, Z => 
                           n5457);
   U2561 : AO4 port map( A => n3775, B => n7334, C => n2416, D => n7326, Z => 
                           n5458);
   U2562 : AO4 port map( A => n3776, B => n7314, C => n2416, D => n7306, Z => 
                           n5459);
   U2563 : AO4 port map( A => n3773, B => n7294, C => n2416, D => n7286, Z => 
                           n5460);
   U2564 : AO4 port map( A => n3774, B => n7274, C => n2416, D => n7266, Z => 
                           n5461);
   U2565 : AO4 port map( A => n3787, B => n7254, C => n2416, D => n7246, Z => 
                           n5462);
   U2566 : AO4 port map( A => n3788, B => n7234, C => n2416, D => n7226, Z => 
                           n5463);
   U2567 : AO4 port map( A => n3785, B => n7214, C => n2416, D => n7206, Z => 
                           n5464);
   U2568 : AO4 port map( A => n3786, B => n7194, C => n2416, D => n7186, Z => 
                           n5465);
   U2569 : AO4 port map( A => n3783, B => n7174, C => n2416, D => n7166, Z => 
                           n5466);
   U2570 : AO4 port map( A => n3784, B => n7154, C => n2416, D => n7146, Z => 
                           n5467);
   U2571 : AO4 port map( A => n3781, B => n7134, C => n2416, D => n7126, Z => 
                           n5468);
   U2572 : AO4 port map( A => n3782, B => n7114, C => n2416, D => n7106, Z => 
                           n5469);
   U2573 : AO4 port map( A => n3795, B => n7094, C => n2416, D => n7086, Z => 
                           n5470);
   U2574 : AO4 port map( A => n3796, B => n7074, C => n2416, D => n7066, Z => 
                           n5471);
   U2575 : AO4 port map( A => n3793, B => n7054, C => n2415, D => n7046, Z => 
                           n5472);
   U2576 : AO4 port map( A => n3794, B => n7034, C => n2415, D => n7026, Z => 
                           n5473);
   U2577 : AO4 port map( A => n3791, B => n7014, C => n2415, D => n7006, Z => 
                           n5474);
   U2578 : AO4 port map( A => n3792, B => n6994, C => n2415, D => n6986, Z => 
                           n5475);
   U2579 : AO4 port map( A => n3789, B => n6974, C => n2415, D => n6966, Z => 
                           n5476);
   U2580 : AO4 port map( A => n3790, B => n6954, C => n2415, D => n6946, Z => 
                           n5477);
   U2581 : AO4 port map( A => n3803, B => n6934, C => n2415, D => n6926, Z => 
                           n5478);
   U2582 : AO4 port map( A => n3804, B => n6914, C => n2415, D => n6906, Z => 
                           n5479);
   U2583 : AO4 port map( A => n3801, B => n6894, C => n2415, D => n6886, Z => 
                           n5480);
   U2584 : AO4 port map( A => n3802, B => n6874, C => n2415, D => n6866, Z => 
                           n5481);
   U2585 : AO4 port map( A => n3799, B => n6854, C => n2415, D => n6846, Z => 
                           n5482);
   U2586 : AO4 port map( A => n3800, B => n6834, C => n2415, D => n6826, Z => 
                           n5483);
   U2587 : AO4 port map( A => n3797, B => n6814, C => n2415, D => n6806, Z => 
                           n5484);
   U2588 : AO4 port map( A => n3798, B => n6794, C => n2415, D => n6786, Z => 
                           n5485);
   U2589 : AO4 port map( A => n3883, B => n7895, C => n2370, D => n7882, Z => 
                           n5942);
   U2590 : AO4 port map( A => n3884, B => n7875, C => n2370, D => n7862, Z => 
                           n5943);
   U2591 : AO4 port map( A => n3881, B => n7855, C => n2370, D => n7842, Z => 
                           n5944);
   U2592 : AO4 port map( A => n3882, B => n7835, C => n2370, D => n7822, Z => 
                           n5945);
   U2593 : AO4 port map( A => n3879, B => n7815, C => n2370, D => n7802, Z => 
                           n5946);
   U2594 : AO4 port map( A => n3880, B => n7795, C => n2370, D => n7782, Z => 
                           n5947);
   U2595 : AO4 port map( A => n3877, B => n7775, C => n2370, D => n7762, Z => 
                           n5948);
   U2596 : AO4 port map( A => n3878, B => n7755, C => n2370, D => n7742, Z => 
                           n5949);
   U2597 : AO4 port map( A => n3891, B => n7735, C => n2370, D => n7722, Z => 
                           n5950);
   U2598 : AO4 port map( A => n3892, B => n7715, C => n2370, D => n7702, Z => 
                           n5951);
   U2599 : AO4 port map( A => n3889, B => n7695, C => n2370, D => n7682, Z => 
                           n5952);
   U2600 : AO4 port map( A => n3890, B => n7675, C => n2370, D => n7662, Z => 
                           n5953);
   U2601 : AO4 port map( A => n3887, B => n7655, C => n2370, D => n7642, Z => 
                           n5954);
   U2602 : AO4 port map( A => n3888, B => n7635, C => n2370, D => n7622, Z => 
                           n5955);
   U2603 : AO4 port map( A => n3885, B => n7615, C => n2369, D => n7602, Z => 
                           n5956);
   U2604 : AO4 port map( A => n3886, B => n7595, C => n2369, D => n7582, Z => 
                           n5957);
   U2605 : AO4 port map( A => n3899, B => n7575, C => n2369, D => n7562, Z => 
                           n5958);
   U2606 : AO4 port map( A => n3900, B => n7555, C => n2369, D => n7542, Z => 
                           n5959);
   U2607 : AO4 port map( A => n3897, B => n7535, C => n2369, D => n7522, Z => 
                           n5960);
   U2608 : AO4 port map( A => n3898, B => n7515, C => n2369, D => n7502, Z => 
                           n5961);
   U2609 : AO4 port map( A => n3895, B => n7495, C => n2369, D => n7482, Z => 
                           n5962);
   U2610 : AO4 port map( A => n3896, B => n7475, C => n2369, D => n7462, Z => 
                           n5963);
   U2611 : AO4 port map( A => n3893, B => n7455, C => n2369, D => n7442, Z => 
                           n5964);
   U2612 : AO4 port map( A => n3894, B => n7435, C => n2369, D => n7422, Z => 
                           n5965);
   U2613 : AO4 port map( A => n3843, B => n7415, C => n2369, D => n7402, Z => 
                           n5966);
   U2614 : AO4 port map( A => n3844, B => n7395, C => n2369, D => n7382, Z => 
                           n5967);
   U2615 : AO4 port map( A => n3841, B => n7375, C => n2369, D => n7362, Z => 
                           n5968);
   U2616 : AO4 port map( A => n3842, B => n7355, C => n2369, D => n7342, Z => 
                           n5969);
   U2617 : AO4 port map( A => n3839, B => n7335, C => n2368, D => n7322, Z => 
                           n5970);
   U2618 : AO4 port map( A => n3840, B => n7315, C => n2368, D => n7302, Z => 
                           n5971);
   U2619 : AO4 port map( A => n3837, B => n7295, C => n2368, D => n7282, Z => 
                           n5972);
   U2620 : AO4 port map( A => n3838, B => n7275, C => n2368, D => n7262, Z => 
                           n5973);
   U2621 : AO4 port map( A => n3851, B => n7255, C => n2368, D => n7242, Z => 
                           n5974);
   U2622 : AO4 port map( A => n3852, B => n7235, C => n2368, D => n7222, Z => 
                           n5975);
   U2623 : AO4 port map( A => n3849, B => n7215, C => n2368, D => n7202, Z => 
                           n5976);
   U2624 : AO4 port map( A => n3850, B => n7195, C => n2368, D => n7182, Z => 
                           n5977);
   U2625 : AO4 port map( A => n3847, B => n7175, C => n2368, D => n7162, Z => 
                           n5978);
   U2626 : AO4 port map( A => n3848, B => n7155, C => n2368, D => n7142, Z => 
                           n5979);
   U2627 : AO4 port map( A => n3845, B => n7135, C => n2368, D => n7122, Z => 
                           n5980);
   U2628 : AO4 port map( A => n3846, B => n7115, C => n2368, D => n7102, Z => 
                           n5981);
   U2629 : AO4 port map( A => n3859, B => n7095, C => n2368, D => n7082, Z => 
                           n5982);
   U2630 : AO4 port map( A => n3860, B => n7075, C => n2368, D => n7062, Z => 
                           n5983);
   U2631 : AO4 port map( A => n3857, B => n7055, C => n2367, D => n7042, Z => 
                           n5984);
   U2632 : AO4 port map( A => n3858, B => n7035, C => n2367, D => n7022, Z => 
                           n5985);
   U2633 : AO4 port map( A => n3855, B => n7015, C => n2367, D => n7002, Z => 
                           n5986);
   U2634 : AO4 port map( A => n3856, B => n6995, C => n2367, D => n6982, Z => 
                           n5987);
   U2635 : AO4 port map( A => n3853, B => n6975, C => n2367, D => n6962, Z => 
                           n5988);
   U2636 : AO4 port map( A => n3854, B => n6955, C => n2367, D => n6942, Z => 
                           n5989);
   U2637 : AO4 port map( A => n3867, B => n6935, C => n2367, D => n6922, Z => 
                           n5990);
   U2638 : AO4 port map( A => n3868, B => n6915, C => n2367, D => n6902, Z => 
                           n5991);
   U2639 : AO4 port map( A => n3865, B => n6895, C => n2367, D => n6882, Z => 
                           n5992);
   U2640 : AO4 port map( A => n3866, B => n6875, C => n2367, D => n6862, Z => 
                           n5993);
   U2641 : AO4 port map( A => n3863, B => n6855, C => n2367, D => n6842, Z => 
                           n5994);
   U2642 : AO4 port map( A => n3864, B => n6835, C => n2367, D => n6822, Z => 
                           n5995);
   U2643 : AO4 port map( A => n3861, B => n6815, C => n2367, D => n6802, Z => 
                           n5996);
   U2644 : AO4 port map( A => n3862, B => n6795, C => n2367, D => n6782, Z => 
                           n5997);
   U2645 : AO4 port map( A => n3947, B => n7896, C => n2322, D => n7878, Z => 
                           n6454);
   U2646 : AO4 port map( A => n3948, B => n7876, C => n2322, D => n7858, Z => 
                           n6455);
   U2647 : AO4 port map( A => n3945, B => n7856, C => n2322, D => n7838, Z => 
                           n6456);
   U2648 : AO4 port map( A => n3946, B => n7836, C => n2322, D => n7818, Z => 
                           n6457);
   U2649 : AO4 port map( A => n3943, B => n7816, C => n2322, D => n7798, Z => 
                           n6458);
   U2650 : AO4 port map( A => n3944, B => n7796, C => n2322, D => n7778, Z => 
                           n6459);
   U2651 : AO4 port map( A => n3941, B => n7776, C => n2322, D => n7758, Z => 
                           n6460);
   U2652 : AO4 port map( A => n3942, B => n7756, C => n2322, D => n7738, Z => 
                           n6461);
   U2653 : AO4 port map( A => n3955, B => n7736, C => n2322, D => n7718, Z => 
                           n6462);
   U2654 : AO4 port map( A => n3956, B => n7716, C => n2322, D => n7698, Z => 
                           n6463);
   U2655 : AO4 port map( A => n3953, B => n7696, C => n2322, D => n7678, Z => 
                           n6464);
   U2656 : AO4 port map( A => n3954, B => n7676, C => n2322, D => n7658, Z => 
                           n6465);
   U2657 : AO4 port map( A => n3951, B => n7656, C => n2322, D => n7638, Z => 
                           n6466);
   U2658 : AO4 port map( A => n3952, B => n7636, C => n2322, D => n7618, Z => 
                           n6467);
   U2659 : AO4 port map( A => n3949, B => n7616, C => n2321, D => n7598, Z => 
                           n6468);
   U2660 : AO4 port map( A => n3950, B => n7596, C => n2321, D => n7578, Z => 
                           n6469);
   U2661 : AO4 port map( A => n3963, B => n7576, C => n2321, D => n7558, Z => 
                           n6470);
   U2662 : AO4 port map( A => n3964, B => n7556, C => n2321, D => n7538, Z => 
                           n6471);
   U2663 : AO4 port map( A => n3961, B => n7536, C => n2321, D => n7518, Z => 
                           n6472);
   U2664 : AO4 port map( A => n3962, B => n7516, C => n2321, D => n7498, Z => 
                           n6473);
   U2665 : AO4 port map( A => n3959, B => n7496, C => n2321, D => n7478, Z => 
                           n6474);
   U2666 : AO4 port map( A => n3960, B => n7476, C => n2321, D => n7458, Z => 
                           n6475);
   U2667 : AO4 port map( A => n3957, B => n7456, C => n2321, D => n7438, Z => 
                           n6476);
   U2668 : AO4 port map( A => n3958, B => n7436, C => n2321, D => n7418, Z => 
                           n6477);
   U2669 : AO4 port map( A => n3907, B => n7416, C => n2321, D => n7398, Z => 
                           n6478);
   U2670 : AO4 port map( A => n3908, B => n7396, C => n2321, D => n7378, Z => 
                           n6479);
   U2671 : AO4 port map( A => n3905, B => n7376, C => n2321, D => n7358, Z => 
                           n6480);
   U2672 : AO4 port map( A => n3906, B => n7356, C => n2321, D => n7338, Z => 
                           n6481);
   U2673 : AO4 port map( A => n3903, B => n7336, C => n2320, D => n7318, Z => 
                           n6482);
   U2674 : AO4 port map( A => n3904, B => n7316, C => n2320, D => n7298, Z => 
                           n6483);
   U2675 : AO4 port map( A => n3901, B => n7296, C => n2320, D => n7278, Z => 
                           n6484);
   U2676 : AO4 port map( A => n3902, B => n7276, C => n2320, D => n7258, Z => 
                           n6485);
   U2677 : AO4 port map( A => n3915, B => n7256, C => n2320, D => n7238, Z => 
                           n6486);
   U2678 : AO4 port map( A => n3916, B => n7236, C => n2320, D => n7218, Z => 
                           n6487);
   U2679 : AO4 port map( A => n3913, B => n7216, C => n2320, D => n7198, Z => 
                           n6488);
   U2680 : AO4 port map( A => n3914, B => n7196, C => n2320, D => n7178, Z => 
                           n6489);
   U2681 : AO4 port map( A => n3911, B => n7176, C => n2320, D => n7158, Z => 
                           n6490);
   U2682 : AO4 port map( A => n3912, B => n7156, C => n2320, D => n7138, Z => 
                           n6491);
   U2683 : AO4 port map( A => n3909, B => n7136, C => n2320, D => n7118, Z => 
                           n6492);
   U2684 : AO4 port map( A => n3910, B => n7116, C => n2320, D => n7098, Z => 
                           n6493);
   U2685 : AO4 port map( A => n3923, B => n7096, C => n2320, D => n7078, Z => 
                           n6494);
   U2686 : AO4 port map( A => n3924, B => n7076, C => n2320, D => n7058, Z => 
                           n6495);
   U2687 : AO4 port map( A => n3921, B => n7056, C => n2319, D => n7038, Z => 
                           n6496);
   U2688 : AO4 port map( A => n3922, B => n7036, C => n2319, D => n7018, Z => 
                           n6497);
   U2689 : AO4 port map( A => n3919, B => n7016, C => n2319, D => n6998, Z => 
                           n6498);
   U2690 : AO4 port map( A => n3920, B => n6996, C => n2319, D => n6978, Z => 
                           n6499);
   U2691 : AO4 port map( A => n3917, B => n6976, C => n2319, D => n6958, Z => 
                           n6500);
   U2692 : AO4 port map( A => n3918, B => n6956, C => n2319, D => n6938, Z => 
                           n6501);
   U2693 : AO4 port map( A => n3931, B => n6936, C => n2319, D => n6918, Z => 
                           n6502);
   U2694 : AO4 port map( A => n3932, B => n6916, C => n2319, D => n6898, Z => 
                           n6503);
   U2695 : AO4 port map( A => n3929, B => n6896, C => n2319, D => n6878, Z => 
                           n6504);
   U2696 : AO4 port map( A => n3930, B => n6876, C => n2319, D => n6858, Z => 
                           n6505);
   U2697 : AO4 port map( A => n3927, B => n6856, C => n2319, D => n6838, Z => 
                           n6506);
   U2698 : AO4 port map( A => n3928, B => n6836, C => n2319, D => n6818, Z => 
                           n6507);
   U2699 : AO4 port map( A => n3925, B => n6816, C => n2319, D => n6798, Z => 
                           n6508);
   U2700 : AO4 port map( A => n3926, B => n6796, C => n2319, D => n6778, Z => 
                           n6509);
   U2701 : AO4 port map( A => n4011, B => n7894, C => n6750, D => n7890, Z => 
                           n4918);
   U2702 : AO4 port map( A => n4012, B => n7874, C => n6750, D => n7870, Z => 
                           n4919);
   U2703 : AO4 port map( A => n4009, B => n7854, C => n6750, D => n7850, Z => 
                           n4920);
   U2704 : AO4 port map( A => n4010, B => n7834, C => n6750, D => n7830, Z => 
                           n4921);
   U2705 : AO4 port map( A => n4007, B => n7814, C => n6750, D => n7810, Z => 
                           n4922);
   U2706 : AO4 port map( A => n4008, B => n7794, C => n6750, D => n7790, Z => 
                           n4923);
   U2707 : AO4 port map( A => n4005, B => n7774, C => n6750, D => n7770, Z => 
                           n4924);
   U2708 : AO4 port map( A => n4006, B => n7754, C => n6750, D => n7750, Z => 
                           n4925);
   U2709 : AO4 port map( A => n4019, B => n7734, C => n6750, D => n7730, Z => 
                           n4926);
   U2710 : AO4 port map( A => n4020, B => n7714, C => n6750, D => n7710, Z => 
                           n4927);
   U2711 : AO4 port map( A => n4017, B => n7694, C => n6750, D => n7690, Z => 
                           n4928);
   U2712 : AO4 port map( A => n4018, B => n7674, C => n6750, D => n7670, Z => 
                           n4929);
   U2713 : AO4 port map( A => n4015, B => n7654, C => n6750, D => n7650, Z => 
                           n4930);
   U2714 : AO4 port map( A => n4016, B => n7634, C => n6750, D => n7630, Z => 
                           n4931);
   U2715 : AO4 port map( A => n4013, B => n7614, C => n6747, D => n7610, Z => 
                           n4932);
   U2716 : AO4 port map( A => n4014, B => n7594, C => n6747, D => n7590, Z => 
                           n4933);
   U2717 : AO4 port map( A => n4027, B => n7574, C => n6747, D => n7570, Z => 
                           n4934);
   U2718 : AO4 port map( A => n4028, B => n7554, C => n6747, D => n7550, Z => 
                           n4935);
   U2719 : AO4 port map( A => n4025, B => n7534, C => n6747, D => n7530, Z => 
                           n4936);
   U2720 : AO4 port map( A => n4026, B => n7514, C => n6747, D => n7510, Z => 
                           n4937);
   U2721 : AO4 port map( A => n4023, B => n7494, C => n6747, D => n7490, Z => 
                           n4938);
   U2722 : AO4 port map( A => n4024, B => n7474, C => n6747, D => n7470, Z => 
                           n4939);
   U2723 : AO4 port map( A => n4021, B => n7454, C => n6747, D => n7450, Z => 
                           n4940);
   U2724 : AO4 port map( A => n4022, B => n7434, C => n6747, D => n7430, Z => 
                           n4941);
   U2725 : AO4 port map( A => n3971, B => n7414, C => n6747, D => n7410, Z => 
                           n4942);
   U2726 : AO4 port map( A => n3972, B => n7394, C => n6747, D => n7390, Z => 
                           n4943);
   U2727 : AO4 port map( A => n3969, B => n7374, C => n6747, D => n7370, Z => 
                           n4944);
   U2728 : AO4 port map( A => n3970, B => n7354, C => n6747, D => n7350, Z => 
                           n4945);
   U2729 : AO4 port map( A => n3967, B => n7334, C => n6746, D => n7330, Z => 
                           n4946);
   U2730 : AO4 port map( A => n3968, B => n7314, C => n6746, D => n7310, Z => 
                           n4947);
   U2731 : AO4 port map( A => n3965, B => n7294, C => n6746, D => n7290, Z => 
                           n4948);
   U2732 : AO4 port map( A => n3966, B => n7274, C => n6746, D => n7270, Z => 
                           n4949);
   U2733 : AO4 port map( A => n3979, B => n7254, C => n6746, D => n7250, Z => 
                           n4950);
   U2734 : AO4 port map( A => n3980, B => n7234, C => n6746, D => n7230, Z => 
                           n4951);
   U2735 : AO4 port map( A => n3977, B => n7214, C => n6746, D => n7210, Z => 
                           n4952);
   U2736 : AO4 port map( A => n3978, B => n7194, C => n6746, D => n7190, Z => 
                           n4953);
   U2737 : AO4 port map( A => n3975, B => n7174, C => n6746, D => n7170, Z => 
                           n4954);
   U2738 : AO4 port map( A => n3976, B => n7154, C => n6746, D => n7150, Z => 
                           n4955);
   U2739 : AO4 port map( A => n3973, B => n7134, C => n6746, D => n7130, Z => 
                           n4956);
   U2740 : AO4 port map( A => n3974, B => n7114, C => n6746, D => n7110, Z => 
                           n4957);
   U2741 : AO4 port map( A => n3987, B => n7094, C => n6746, D => n7090, Z => 
                           n4958);
   U2742 : AO4 port map( A => n3988, B => n7074, C => n6746, D => n7070, Z => 
                           n4959);
   U2743 : AO4 port map( A => n3985, B => n7054, C => n6745, D => n7050, Z => 
                           n4960);
   U2744 : AO4 port map( A => n3986, B => n7034, C => n6745, D => n7030, Z => 
                           n4961);
   U2745 : AO4 port map( A => n3983, B => n7014, C => n6745, D => n7010, Z => 
                           n4962);
   U2746 : AO4 port map( A => n3984, B => n6994, C => n6745, D => n6990, Z => 
                           n4963);
   U2747 : AO4 port map( A => n3981, B => n6974, C => n6745, D => n6970, Z => 
                           n4964);
   U2748 : AO4 port map( A => n3982, B => n6954, C => n6745, D => n6950, Z => 
                           n4965);
   U2749 : AO4 port map( A => n3995, B => n6934, C => n6745, D => n6930, Z => 
                           n4966);
   U2750 : AO4 port map( A => n3996, B => n6914, C => n6745, D => n6910, Z => 
                           n4967);
   U2751 : AO4 port map( A => n3993, B => n6894, C => n6745, D => n6890, Z => 
                           n4968);
   U2752 : AO4 port map( A => n3994, B => n6874, C => n6745, D => n6870, Z => 
                           n4969);
   U2753 : AO4 port map( A => n3991, B => n6854, C => n6745, D => n6850, Z => 
                           n4970);
   U2754 : AO4 port map( A => n3992, B => n6834, C => n6745, D => n6830, Z => 
                           n4971);
   U2755 : AO4 port map( A => n3989, B => n6814, C => n6745, D => n6810, Z => 
                           n4972);
   U2756 : AO4 port map( A => n3990, B => n6794, C => n6745, D => n6790, Z => 
                           n4973);
   U2757 : AO4 port map( A => n4075, B => n7895, C => n2412, D => n7885, Z => 
                           n5494);
   U2758 : AO4 port map( A => n4076, B => n7875, C => n2412, D => n7865, Z => 
                           n5495);
   U2759 : AO4 port map( A => n4073, B => n7855, C => n2412, D => n7845, Z => 
                           n5496);
   U2760 : AO4 port map( A => n4074, B => n7835, C => n2412, D => n7825, Z => 
                           n5497);
   U2761 : AO4 port map( A => n4071, B => n7815, C => n2412, D => n7805, Z => 
                           n5498);
   U2762 : AO4 port map( A => n4072, B => n7795, C => n2412, D => n7785, Z => 
                           n5499);
   U2763 : AO4 port map( A => n4069, B => n7775, C => n2412, D => n7765, Z => 
                           n5500);
   U2764 : AO4 port map( A => n4070, B => n7755, C => n2412, D => n7745, Z => 
                           n5501);
   U2765 : AO4 port map( A => n4083, B => n7735, C => n2412, D => n7725, Z => 
                           n5502);
   U2766 : AO4 port map( A => n4084, B => n7715, C => n2412, D => n7705, Z => 
                           n5503);
   U2767 : AO4 port map( A => n4081, B => n7695, C => n2412, D => n7685, Z => 
                           n5504);
   U2768 : AO4 port map( A => n4082, B => n7675, C => n2412, D => n7665, Z => 
                           n5505);
   U2769 : AO4 port map( A => n4079, B => n7655, C => n2412, D => n7645, Z => 
                           n5506);
   U2770 : AO4 port map( A => n4080, B => n7635, C => n2412, D => n7625, Z => 
                           n5507);
   U2771 : AO4 port map( A => n4077, B => n7615, C => n2411, D => n7605, Z => 
                           n5508);
   U2772 : AO4 port map( A => n4078, B => n7595, C => n2411, D => n7585, Z => 
                           n5509);
   U2773 : AO4 port map( A => n4091, B => n7575, C => n2411, D => n7565, Z => 
                           n5510);
   U2774 : AO4 port map( A => n4092, B => n7555, C => n2411, D => n7545, Z => 
                           n5511);
   U2775 : AO4 port map( A => n4089, B => n7535, C => n2411, D => n7525, Z => 
                           n5512);
   U2776 : AO4 port map( A => n4090, B => n7515, C => n2411, D => n7505, Z => 
                           n5513);
   U2777 : AO4 port map( A => n4087, B => n7495, C => n2411, D => n7485, Z => 
                           n5514);
   U2778 : AO4 port map( A => n4088, B => n7475, C => n2411, D => n7465, Z => 
                           n5515);
   U2779 : AO4 port map( A => n4085, B => n7455, C => n2411, D => n7445, Z => 
                           n5516);
   U2780 : AO4 port map( A => n4086, B => n7435, C => n2411, D => n7425, Z => 
                           n5517);
   U2781 : AO4 port map( A => n4035, B => n7415, C => n2411, D => n7405, Z => 
                           n5518);
   U2782 : AO4 port map( A => n4036, B => n7395, C => n2411, D => n7385, Z => 
                           n5519);
   U2783 : AO4 port map( A => n4033, B => n7375, C => n2411, D => n7365, Z => 
                           n5520);
   U2784 : AO4 port map( A => n4034, B => n7355, C => n2411, D => n7345, Z => 
                           n5521);
   U2785 : AO4 port map( A => n4031, B => n7335, C => n2410, D => n7325, Z => 
                           n5522);
   U2786 : AO4 port map( A => n4032, B => n7315, C => n2410, D => n7305, Z => 
                           n5523);
   U2787 : AO4 port map( A => n4029, B => n7295, C => n2410, D => n7285, Z => 
                           n5524);
   U2788 : AO4 port map( A => n4030, B => n7275, C => n2410, D => n7265, Z => 
                           n5525);
   U2789 : AO4 port map( A => n4043, B => n7255, C => n2410, D => n7245, Z => 
                           n5526);
   U2790 : AO4 port map( A => n4044, B => n7235, C => n2410, D => n7225, Z => 
                           n5527);
   U2791 : AO4 port map( A => n4041, B => n7215, C => n2410, D => n7205, Z => 
                           n5528);
   U2792 : AO4 port map( A => n4042, B => n7195, C => n2410, D => n7185, Z => 
                           n5529);
   U2793 : AO4 port map( A => n4039, B => n7175, C => n2410, D => n7165, Z => 
                           n5530);
   U2794 : AO4 port map( A => n4040, B => n7155, C => n2410, D => n7145, Z => 
                           n5531);
   U2795 : AO4 port map( A => n4037, B => n7135, C => n2410, D => n7125, Z => 
                           n5532);
   U2796 : AO4 port map( A => n4038, B => n7115, C => n2410, D => n7105, Z => 
                           n5533);
   U2797 : AO4 port map( A => n4051, B => n7095, C => n2410, D => n7085, Z => 
                           n5534);
   U2798 : AO4 port map( A => n4052, B => n7075, C => n2410, D => n7065, Z => 
                           n5535);
   U2799 : AO4 port map( A => n4049, B => n7055, C => n2409, D => n7045, Z => 
                           n5536);
   U2800 : AO4 port map( A => n4050, B => n7035, C => n2409, D => n7025, Z => 
                           n5537);
   U2801 : AO4 port map( A => n4047, B => n7015, C => n2409, D => n7005, Z => 
                           n5538);
   U2802 : AO4 port map( A => n4048, B => n6995, C => n2409, D => n6985, Z => 
                           n5539);
   U2803 : AO4 port map( A => n4045, B => n6975, C => n2409, D => n6965, Z => 
                           n5540);
   U2804 : AO4 port map( A => n4046, B => n6955, C => n2409, D => n6945, Z => 
                           n5541);
   U2805 : AO4 port map( A => n4059, B => n6935, C => n2409, D => n6925, Z => 
                           n5542);
   U2806 : AO4 port map( A => n4060, B => n6915, C => n2409, D => n6905, Z => 
                           n5543);
   U2807 : AO4 port map( A => n4057, B => n6895, C => n2409, D => n6885, Z => 
                           n5544);
   U2808 : AO4 port map( A => n4058, B => n6875, C => n2409, D => n6865, Z => 
                           n5545);
   U2809 : AO4 port map( A => n4055, B => n6855, C => n2409, D => n6845, Z => 
                           n5546);
   U2810 : AO4 port map( A => n4056, B => n6835, C => n2409, D => n6825, Z => 
                           n5547);
   U2811 : AO4 port map( A => n4053, B => n6815, C => n2409, D => n6805, Z => 
                           n5548);
   U2812 : AO4 port map( A => n4054, B => n6795, C => n2409, D => n6785, Z => 
                           n5549);
   U2813 : AO4 port map( A => n4139, B => n7895, C => n2364, D => n7881, Z => 
                           n6006);
   U2814 : AO4 port map( A => n4140, B => n7875, C => n2364, D => n7861, Z => 
                           n6007);
   U2815 : AO4 port map( A => n4137, B => n7855, C => n2364, D => n7841, Z => 
                           n6008);
   U2816 : AO4 port map( A => n4138, B => n7835, C => n2364, D => n7821, Z => 
                           n6009);
   U2817 : AO4 port map( A => n4135, B => n7815, C => n2364, D => n7801, Z => 
                           n6010);
   U2818 : AO4 port map( A => n4136, B => n7795, C => n2364, D => n7781, Z => 
                           n6011);
   U2819 : AO4 port map( A => n4133, B => n7775, C => n2364, D => n7761, Z => 
                           n6012);
   U2820 : AO4 port map( A => n4134, B => n7755, C => n2364, D => n7741, Z => 
                           n6013);
   U2821 : AO4 port map( A => n4147, B => n7735, C => n2364, D => n7721, Z => 
                           n6014);
   U2822 : AO4 port map( A => n4148, B => n7715, C => n2364, D => n7701, Z => 
                           n6015);
   U2823 : AO4 port map( A => n4145, B => n7695, C => n2364, D => n7681, Z => 
                           n6016);
   U2824 : AO4 port map( A => n4146, B => n7675, C => n2364, D => n7661, Z => 
                           n6017);
   U2825 : AO4 port map( A => n4143, B => n7655, C => n2364, D => n7641, Z => 
                           n6018);
   U2826 : AO4 port map( A => n4144, B => n7635, C => n2364, D => n7621, Z => 
                           n6019);
   U2827 : AO4 port map( A => n4141, B => n7615, C => n2363, D => n7601, Z => 
                           n6020);
   U2828 : AO4 port map( A => n4142, B => n7595, C => n2363, D => n7581, Z => 
                           n6021);
   U2829 : AO4 port map( A => n4155, B => n7575, C => n2363, D => n7561, Z => 
                           n6022);
   U2830 : AO4 port map( A => n4156, B => n7555, C => n2363, D => n7541, Z => 
                           n6023);
   U2831 : AO4 port map( A => n4153, B => n7535, C => n2363, D => n7521, Z => 
                           n6024);
   U2832 : AO4 port map( A => n4154, B => n7515, C => n2363, D => n7501, Z => 
                           n6025);
   U2833 : AO4 port map( A => n4151, B => n7495, C => n2363, D => n7481, Z => 
                           n6026);
   U2834 : AO4 port map( A => n4152, B => n7475, C => n2363, D => n7461, Z => 
                           n6027);
   U2835 : AO4 port map( A => n4149, B => n7455, C => n2363, D => n7441, Z => 
                           n6028);
   U2836 : AO4 port map( A => n4150, B => n7435, C => n2363, D => n7421, Z => 
                           n6029);
   U2837 : AO4 port map( A => n4099, B => n7415, C => n2363, D => n7401, Z => 
                           n6030);
   U2838 : AO4 port map( A => n4100, B => n7395, C => n2363, D => n7381, Z => 
                           n6031);
   U2839 : AO4 port map( A => n4097, B => n7375, C => n2363, D => n7361, Z => 
                           n6032);
   U2840 : AO4 port map( A => n4098, B => n7355, C => n2363, D => n7341, Z => 
                           n6033);
   U2841 : AO4 port map( A => n4095, B => n7335, C => n2362, D => n7321, Z => 
                           n6034);
   U2842 : AO4 port map( A => n4096, B => n7315, C => n2362, D => n7301, Z => 
                           n6035);
   U2843 : AO4 port map( A => n4093, B => n7295, C => n2362, D => n7281, Z => 
                           n6036);
   U2844 : AO4 port map( A => n4094, B => n7275, C => n2362, D => n7261, Z => 
                           n6037);
   U2845 : AO4 port map( A => n4107, B => n7255, C => n2362, D => n7241, Z => 
                           n6038);
   U2846 : AO4 port map( A => n4108, B => n7235, C => n2362, D => n7221, Z => 
                           n6039);
   U2847 : AO4 port map( A => n4105, B => n7215, C => n2362, D => n7201, Z => 
                           n6040);
   U2848 : AO4 port map( A => n4106, B => n7195, C => n2362, D => n7181, Z => 
                           n6041);
   U2849 : AO4 port map( A => n4103, B => n7175, C => n2362, D => n7161, Z => 
                           n6042);
   U2850 : AO4 port map( A => n4104, B => n7155, C => n2362, D => n7141, Z => 
                           n6043);
   U2851 : AO4 port map( A => n4101, B => n7135, C => n2362, D => n7121, Z => 
                           n6044);
   U2852 : AO4 port map( A => n4102, B => n7115, C => n2362, D => n7101, Z => 
                           n6045);
   U2853 : AO4 port map( A => n4115, B => n7095, C => n2362, D => n7081, Z => 
                           n6046);
   U2854 : AO4 port map( A => n4116, B => n7075, C => n2362, D => n7061, Z => 
                           n6047);
   U2855 : AO4 port map( A => n4113, B => n7055, C => n2361, D => n7041, Z => 
                           n6048);
   U2856 : AO4 port map( A => n4114, B => n7035, C => n2361, D => n7021, Z => 
                           n6049);
   U2857 : AO4 port map( A => n4111, B => n7015, C => n2361, D => n7001, Z => 
                           n6050);
   U2858 : AO4 port map( A => n4112, B => n6995, C => n2361, D => n6981, Z => 
                           n6051);
   U2859 : AO4 port map( A => n4109, B => n6975, C => n2361, D => n6961, Z => 
                           n6052);
   U2860 : AO4 port map( A => n4110, B => n6955, C => n2361, D => n6941, Z => 
                           n6053);
   U2861 : AO4 port map( A => n4123, B => n6935, C => n2361, D => n6921, Z => 
                           n6054);
   U2862 : AO4 port map( A => n4124, B => n6915, C => n2361, D => n6901, Z => 
                           n6055);
   U2863 : AO4 port map( A => n4121, B => n6895, C => n2361, D => n6881, Z => 
                           n6056);
   U2864 : AO4 port map( A => n4122, B => n6875, C => n2361, D => n6861, Z => 
                           n6057);
   U2865 : AO4 port map( A => n4119, B => n6855, C => n2361, D => n6841, Z => 
                           n6058);
   U2866 : AO4 port map( A => n4120, B => n6835, C => n2361, D => n6821, Z => 
                           n6059);
   U2867 : AO4 port map( A => n4117, B => n6815, C => n2361, D => n6801, Z => 
                           n6060);
   U2868 : AO4 port map( A => n4118, B => n6795, C => n2361, D => n6781, Z => 
                           n6061);
   U2869 : AO4 port map( A => n4203, B => n7896, C => n2316, D => n7877, Z => 
                           n6518);
   U2870 : AO4 port map( A => n4204, B => n7876, C => n2316, D => n7857, Z => 
                           n6519);
   U2871 : AO4 port map( A => n4201, B => n7856, C => n2316, D => n7837, Z => 
                           n6520);
   U2872 : AO4 port map( A => n4202, B => n7836, C => n2316, D => n7817, Z => 
                           n6521);
   U2873 : AO4 port map( A => n4199, B => n7816, C => n2316, D => n7797, Z => 
                           n6522);
   U2874 : AO4 port map( A => n4200, B => n7796, C => n2316, D => n7777, Z => 
                           n6523);
   U2875 : AO4 port map( A => n4197, B => n7776, C => n2316, D => n7757, Z => 
                           n6524);
   U2876 : AO4 port map( A => n4198, B => n7756, C => n2316, D => n7737, Z => 
                           n6525);
   U2877 : AO4 port map( A => n4211, B => n7736, C => n2316, D => n7717, Z => 
                           n6526);
   U2878 : AO4 port map( A => n4212, B => n7716, C => n2316, D => n7697, Z => 
                           n6527);
   U2879 : AO4 port map( A => n4209, B => n7696, C => n2316, D => n7677, Z => 
                           n6528);
   U2880 : AO4 port map( A => n4210, B => n7676, C => n2316, D => n7657, Z => 
                           n6529);
   U2881 : AO4 port map( A => n4207, B => n7656, C => n2316, D => n7637, Z => 
                           n6530);
   U2882 : AO4 port map( A => n4208, B => n7636, C => n2316, D => n7617, Z => 
                           n6531);
   U2883 : AO4 port map( A => n4205, B => n7616, C => n2315, D => n7597, Z => 
                           n6532);
   U2884 : AO4 port map( A => n4206, B => n7596, C => n2315, D => n7577, Z => 
                           n6533);
   U2885 : AO4 port map( A => n4219, B => n7576, C => n2315, D => n7557, Z => 
                           n6534);
   U2886 : AO4 port map( A => n4220, B => n7556, C => n2315, D => n7537, Z => 
                           n6535);
   U2887 : AO4 port map( A => n4217, B => n7536, C => n2315, D => n7517, Z => 
                           n6536);
   U2888 : AO4 port map( A => n4218, B => n7516, C => n2315, D => n7497, Z => 
                           n6537);
   U2889 : AO4 port map( A => n4215, B => n7496, C => n2315, D => n7477, Z => 
                           n6538);
   U2890 : AO4 port map( A => n4216, B => n7476, C => n2315, D => n7457, Z => 
                           n6539);
   U2891 : AO4 port map( A => n4213, B => n7456, C => n2315, D => n7437, Z => 
                           n6540);
   U2892 : AO4 port map( A => n4214, B => n7436, C => n2315, D => n7417, Z => 
                           n6541);
   U2893 : AO4 port map( A => n4163, B => n7416, C => n2315, D => n7397, Z => 
                           n6542);
   U2894 : AO4 port map( A => n4164, B => n7396, C => n2315, D => n7377, Z => 
                           n6543);
   U2895 : AO4 port map( A => n4161, B => n7376, C => n2315, D => n7357, Z => 
                           n6544);
   U2896 : AO4 port map( A => n4162, B => n7356, C => n2315, D => n7337, Z => 
                           n6545);
   U2897 : AO4 port map( A => n4159, B => n7336, C => n2314, D => n7317, Z => 
                           n6546);
   U2898 : AO4 port map( A => n4160, B => n7316, C => n2314, D => n7297, Z => 
                           n6547);
   U2899 : AO4 port map( A => n4157, B => n7296, C => n2314, D => n7277, Z => 
                           n6548);
   U2900 : AO4 port map( A => n4158, B => n7276, C => n2314, D => n7257, Z => 
                           n6549);
   U2901 : AO4 port map( A => n4171, B => n7256, C => n2314, D => n7237, Z => 
                           n6550);
   U2902 : AO4 port map( A => n4172, B => n7236, C => n2314, D => n7217, Z => 
                           n6551);
   U2903 : AO4 port map( A => n4169, B => n7216, C => n2314, D => n7197, Z => 
                           n6552);
   U2904 : AO4 port map( A => n4170, B => n7196, C => n2314, D => n7177, Z => 
                           n6553);
   U2905 : AO4 port map( A => n4167, B => n7176, C => n2314, D => n7157, Z => 
                           n6554);
   U2906 : AO4 port map( A => n4168, B => n7156, C => n2314, D => n7137, Z => 
                           n6555);
   U2907 : AO4 port map( A => n4165, B => n7136, C => n2314, D => n7117, Z => 
                           n6556);
   U2908 : AO4 port map( A => n4166, B => n7116, C => n2314, D => n7097, Z => 
                           n6557);
   U2909 : AO4 port map( A => n4179, B => n7096, C => n2314, D => n7077, Z => 
                           n6558);
   U2910 : AO4 port map( A => n4180, B => n7076, C => n2314, D => n7057, Z => 
                           n6559);
   U2911 : AO4 port map( A => n4177, B => n7056, C => n2313, D => n7037, Z => 
                           n6560);
   U2912 : AO4 port map( A => n4178, B => n7036, C => n2313, D => n7017, Z => 
                           n6561);
   U2913 : AO4 port map( A => n4175, B => n7016, C => n2313, D => n6997, Z => 
                           n6562);
   U2914 : AO4 port map( A => n4176, B => n6996, C => n2313, D => n6977, Z => 
                           n6563);
   U2915 : AO4 port map( A => n4173, B => n6976, C => n2313, D => n6957, Z => 
                           n6564);
   U2916 : AO4 port map( A => n4174, B => n6956, C => n2313, D => n6937, Z => 
                           n6565);
   U2917 : AO4 port map( A => n4187, B => n6936, C => n2313, D => n6917, Z => 
                           n6566);
   U2918 : AO4 port map( A => n4188, B => n6916, C => n2313, D => n6897, Z => 
                           n6567);
   U2919 : AO4 port map( A => n4185, B => n6896, C => n2313, D => n6877, Z => 
                           n6568);
   U2920 : AO4 port map( A => n4186, B => n6876, C => n2313, D => n6857, Z => 
                           n6569);
   U2921 : AO4 port map( A => n4183, B => n6856, C => n2313, D => n6837, Z => 
                           n6570);
   U2922 : AO4 port map( A => n4184, B => n6836, C => n2313, D => n6817, Z => 
                           n6571);
   U2923 : AO4 port map( A => n4181, B => n6816, C => n2313, D => n6797, Z => 
                           n6572);
   U2924 : AO4 port map( A => n4182, B => n6796, C => n2313, D => n6777, Z => 
                           n6573);
   U2925 : AO4 port map( A => n4267, B => n7894, C => n6742, D => n7889, Z => 
                           n4982);
   U2926 : AO4 port map( A => n4268, B => n7874, C => n6742, D => n7869, Z => 
                           n4983);
   U2927 : AO4 port map( A => n4265, B => n7854, C => n6742, D => n7849, Z => 
                           n4984);
   U2928 : AO4 port map( A => n4266, B => n7834, C => n6742, D => n7829, Z => 
                           n4985);
   U2929 : AO4 port map( A => n4263, B => n7814, C => n6742, D => n7809, Z => 
                           n4986);
   U2930 : AO4 port map( A => n4264, B => n7794, C => n6742, D => n7789, Z => 
                           n4987);
   U2931 : AO4 port map( A => n4261, B => n7774, C => n6742, D => n7769, Z => 
                           n4988);
   U2932 : AO4 port map( A => n4262, B => n7754, C => n6742, D => n7749, Z => 
                           n4989);
   U2933 : AO4 port map( A => n4275, B => n7734, C => n6742, D => n7729, Z => 
                           n4990);
   U2934 : AO4 port map( A => n4276, B => n7714, C => n6742, D => n7709, Z => 
                           n4991);
   U2935 : AO4 port map( A => n4273, B => n7694, C => n6742, D => n7689, Z => 
                           n4992);
   U2936 : AO4 port map( A => n4274, B => n7674, C => n6742, D => n7669, Z => 
                           n4993);
   U2937 : AO4 port map( A => n4271, B => n7654, C => n6742, D => n7649, Z => 
                           n4994);
   U2938 : AO4 port map( A => n4272, B => n7634, C => n6742, D => n7629, Z => 
                           n4995);
   U2939 : AO4 port map( A => n4269, B => n7614, C => n6741, D => n7609, Z => 
                           n4996);
   U2940 : AO4 port map( A => n4270, B => n7594, C => n6741, D => n7589, Z => 
                           n4997);
   U2941 : AO4 port map( A => n4283, B => n7574, C => n6741, D => n7569, Z => 
                           n4998);
   U2942 : AO4 port map( A => n4284, B => n7554, C => n6741, D => n7549, Z => 
                           n4999);
   U2943 : AO4 port map( A => n4281, B => n7534, C => n6741, D => n7529, Z => 
                           n5000);
   U2944 : AO4 port map( A => n4282, B => n7514, C => n6741, D => n7509, Z => 
                           n5001);
   U2945 : AO4 port map( A => n4279, B => n7494, C => n6741, D => n7489, Z => 
                           n5002);
   U2946 : AO4 port map( A => n4280, B => n7474, C => n6741, D => n7469, Z => 
                           n5003);
   U2947 : AO4 port map( A => n4277, B => n7454, C => n6741, D => n7449, Z => 
                           n5004);
   U2948 : AO4 port map( A => n4278, B => n7434, C => n6741, D => n7429, Z => 
                           n5005);
   U2949 : AO4 port map( A => n4227, B => n7414, C => n6741, D => n7409, Z => 
                           n5006);
   U2950 : AO4 port map( A => n4228, B => n7394, C => n6741, D => n7389, Z => 
                           n5007);
   U2951 : AO4 port map( A => n4225, B => n7374, C => n6741, D => n7369, Z => 
                           n5008);
   U2952 : AO4 port map( A => n4226, B => n7354, C => n6741, D => n7349, Z => 
                           n5009);
   U2953 : AO4 port map( A => n4223, B => n7334, C => n6740, D => n7329, Z => 
                           n5010);
   U2954 : AO4 port map( A => n4224, B => n7314, C => n6740, D => n7309, Z => 
                           n5011);
   U2955 : AO4 port map( A => n4221, B => n7294, C => n6740, D => n7289, Z => 
                           n5012);
   U2956 : AO4 port map( A => n4222, B => n7274, C => n6740, D => n7269, Z => 
                           n5013);
   U2957 : AO4 port map( A => n4235, B => n7254, C => n6740, D => n7249, Z => 
                           n5014);
   U2958 : AO4 port map( A => n4236, B => n7234, C => n6740, D => n7229, Z => 
                           n5015);
   U2959 : AO4 port map( A => n4233, B => n7214, C => n6740, D => n7209, Z => 
                           n5016);
   U2960 : AO4 port map( A => n4234, B => n7194, C => n6740, D => n7189, Z => 
                           n5017);
   U2961 : AO4 port map( A => n4231, B => n7174, C => n6740, D => n7169, Z => 
                           n5018);
   U2962 : AO4 port map( A => n4232, B => n7154, C => n6740, D => n7149, Z => 
                           n5019);
   U2963 : AO4 port map( A => n4229, B => n7134, C => n6740, D => n7129, Z => 
                           n5020);
   U2964 : AO4 port map( A => n4230, B => n7114, C => n6740, D => n7109, Z => 
                           n5021);
   U2965 : AO4 port map( A => n4243, B => n7094, C => n6740, D => n7089, Z => 
                           n5022);
   U2966 : AO4 port map( A => n4244, B => n7074, C => n6740, D => n7069, Z => 
                           n5023);
   U2967 : AO4 port map( A => n4241, B => n7054, C => n6739, D => n7049, Z => 
                           n5024);
   U2968 : AO4 port map( A => n4242, B => n7034, C => n6739, D => n7029, Z => 
                           n5025);
   U2969 : AO4 port map( A => n4239, B => n7014, C => n6739, D => n7009, Z => 
                           n5026);
   U2970 : AO4 port map( A => n4240, B => n6994, C => n6739, D => n6989, Z => 
                           n5027);
   U2971 : AO4 port map( A => n4237, B => n6974, C => n6739, D => n6969, Z => 
                           n5028);
   U2972 : AO4 port map( A => n4238, B => n6954, C => n6739, D => n6949, Z => 
                           n5029);
   U2973 : AO4 port map( A => n4251, B => n6934, C => n6739, D => n6929, Z => 
                           n5030);
   U2974 : AO4 port map( A => n4252, B => n6914, C => n6739, D => n6909, Z => 
                           n5031);
   U2975 : AO4 port map( A => n4249, B => n6894, C => n6739, D => n6889, Z => 
                           n5032);
   U2976 : AO4 port map( A => n4250, B => n6874, C => n6739, D => n6869, Z => 
                           n5033);
   U2977 : AO4 port map( A => n4247, B => n6854, C => n6739, D => n6849, Z => 
                           n5034);
   U2978 : AO4 port map( A => n4248, B => n6834, C => n6739, D => n6829, Z => 
                           n5035);
   U2979 : AO4 port map( A => n4245, B => n6814, C => n6739, D => n6809, Z => 
                           n5036);
   U2980 : AO4 port map( A => n4246, B => n6794, C => n6739, D => n6789, Z => 
                           n5037);
   U2981 : AO4 port map( A => n4332, B => n7895, C => n2406, D => n7885, Z => 
                           n5558);
   U2982 : AO4 port map( A => n4333, B => n7875, C => n2406, D => n7865, Z => 
                           n5559);
   U2983 : AO4 port map( A => n4330, B => n7855, C => n2406, D => n7845, Z => 
                           n5560);
   U2984 : AO4 port map( A => n4331, B => n7835, C => n2406, D => n7825, Z => 
                           n5561);
   U2985 : AO4 port map( A => n4328, B => n7815, C => n2406, D => n7805, Z => 
                           n5562);
   U2986 : AO4 port map( A => n4329, B => n7795, C => n2406, D => n7785, Z => 
                           n5563);
   U2987 : AO4 port map( A => n4326, B => n7775, C => n2406, D => n7765, Z => 
                           n5564);
   U2988 : AO4 port map( A => n4327, B => n7755, C => n2406, D => n7745, Z => 
                           n5565);
   U2989 : AO4 port map( A => n4340, B => n7735, C => n2406, D => n7725, Z => 
                           n5566);
   U2990 : AO4 port map( A => n4341, B => n7715, C => n2406, D => n7705, Z => 
                           n5567);
   U2991 : AO4 port map( A => n4338, B => n7695, C => n2406, D => n7685, Z => 
                           n5568);
   U2992 : AO4 port map( A => n4339, B => n7675, C => n2406, D => n7665, Z => 
                           n5569);
   U2993 : AO4 port map( A => n4336, B => n7655, C => n2406, D => n7645, Z => 
                           n5570);
   U2994 : AO4 port map( A => n4337, B => n7635, C => n2406, D => n7625, Z => 
                           n5571);
   U2995 : AO4 port map( A => n4334, B => n7615, C => n2405, D => n7605, Z => 
                           n5572);
   U2996 : AO4 port map( A => n4335, B => n7595, C => n2405, D => n7585, Z => 
                           n5573);
   U2997 : AO4 port map( A => n4348, B => n7575, C => n2405, D => n7565, Z => 
                           n5574);
   U2998 : AO4 port map( A => n4349, B => n7555, C => n2405, D => n7545, Z => 
                           n5575);
   U2999 : AO4 port map( A => n4346, B => n7535, C => n2405, D => n7525, Z => 
                           n5576);
   U3000 : AO4 port map( A => n4347, B => n7515, C => n2405, D => n7505, Z => 
                           n5577);
   U3001 : AO4 port map( A => n4344, B => n7495, C => n2405, D => n7485, Z => 
                           n5578);
   U3002 : AO4 port map( A => n4345, B => n7475, C => n2405, D => n7465, Z => 
                           n5579);
   U3003 : AO4 port map( A => n4342, B => n7455, C => n2405, D => n7445, Z => 
                           n5580);
   U3004 : AO4 port map( A => n4343, B => n7435, C => n2405, D => n7425, Z => 
                           n5581);
   U3005 : AO4 port map( A => n4292, B => n7415, C => n2405, D => n7405, Z => 
                           n5582);
   U3006 : AO4 port map( A => n4293, B => n7395, C => n2405, D => n7385, Z => 
                           n5583);
   U3007 : AO4 port map( A => n4290, B => n7375, C => n2405, D => n7365, Z => 
                           n5584);
   U3008 : AO4 port map( A => n4291, B => n7355, C => n2405, D => n7345, Z => 
                           n5585);
   U3009 : AO4 port map( A => n4288, B => n7335, C => n2404, D => n7325, Z => 
                           n5586);
   U3010 : AO4 port map( A => n4289, B => n7315, C => n2404, D => n7305, Z => 
                           n5587);
   U3011 : AO4 port map( A => n4286, B => n7295, C => n2404, D => n7285, Z => 
                           n5588);
   U3012 : AO4 port map( A => n4287, B => n7275, C => n2404, D => n7265, Z => 
                           n5589);
   U3013 : AO4 port map( A => n4300, B => n7255, C => n2404, D => n7245, Z => 
                           n5590);
   U3014 : AO4 port map( A => n4301, B => n7235, C => n2404, D => n7225, Z => 
                           n5591);
   U3015 : AO4 port map( A => n4298, B => n7215, C => n2404, D => n7205, Z => 
                           n5592);
   U3016 : AO4 port map( A => n4299, B => n7195, C => n2404, D => n7185, Z => 
                           n5593);
   U3017 : AO4 port map( A => n4296, B => n7175, C => n2404, D => n7165, Z => 
                           n5594);
   U3018 : AO4 port map( A => n4297, B => n7155, C => n2404, D => n7145, Z => 
                           n5595);
   U3019 : AO4 port map( A => n4294, B => n7135, C => n2404, D => n7125, Z => 
                           n5596);
   U3020 : AO4 port map( A => n4295, B => n7115, C => n2404, D => n7105, Z => 
                           n5597);
   U3021 : AO4 port map( A => n4308, B => n7095, C => n2404, D => n7085, Z => 
                           n5598);
   U3022 : AO4 port map( A => n4309, B => n7075, C => n2404, D => n7065, Z => 
                           n5599);
   U3023 : AO4 port map( A => n4306, B => n7055, C => n2403, D => n7045, Z => 
                           n5600);
   U3024 : AO4 port map( A => n4307, B => n7035, C => n2403, D => n7025, Z => 
                           n5601);
   U3025 : AO4 port map( A => n4304, B => n7015, C => n2403, D => n7005, Z => 
                           n5602);
   U3026 : AO4 port map( A => n4305, B => n6995, C => n2403, D => n6985, Z => 
                           n5603);
   U3027 : AO4 port map( A => n4302, B => n6975, C => n2403, D => n6965, Z => 
                           n5604);
   U3028 : AO4 port map( A => n4303, B => n6955, C => n2403, D => n6945, Z => 
                           n5605);
   U3029 : AO4 port map( A => n4316, B => n6935, C => n2403, D => n6925, Z => 
                           n5606);
   U3030 : AO4 port map( A => n4317, B => n6915, C => n2403, D => n6905, Z => 
                           n5607);
   U3031 : AO4 port map( A => n4314, B => n6895, C => n2403, D => n6885, Z => 
                           n5608);
   U3032 : AO4 port map( A => n4315, B => n6875, C => n2403, D => n6865, Z => 
                           n5609);
   U3033 : AO4 port map( A => n4312, B => n6855, C => n2403, D => n6845, Z => 
                           n5610);
   U3034 : AO4 port map( A => n4313, B => n6835, C => n2403, D => n6825, Z => 
                           n5611);
   U3035 : AO4 port map( A => n4310, B => n6815, C => n2403, D => n6805, Z => 
                           n5612);
   U3036 : AO4 port map( A => n4311, B => n6795, C => n2403, D => n6785, Z => 
                           n5613);
   U3037 : AO4 port map( A => n4396, B => n7895, C => n2358, D => n7881, Z => 
                           n6070);
   U3038 : AO4 port map( A => n4397, B => n7875, C => n2358, D => n7861, Z => 
                           n6071);
   U3039 : AO4 port map( A => n4394, B => n7855, C => n2358, D => n7841, Z => 
                           n6072);
   U3040 : AO4 port map( A => n4395, B => n7835, C => n2358, D => n7821, Z => 
                           n6073);
   U3041 : AO4 port map( A => n4392, B => n7815, C => n2358, D => n7801, Z => 
                           n6074);
   U3042 : AO4 port map( A => n4393, B => n7795, C => n2358, D => n7781, Z => 
                           n6075);
   U3043 : AO4 port map( A => n4390, B => n7775, C => n2358, D => n7761, Z => 
                           n6076);
   U3044 : AO4 port map( A => n4391, B => n7755, C => n2358, D => n7741, Z => 
                           n6077);
   U3045 : AO4 port map( A => n4404, B => n7735, C => n2358, D => n7721, Z => 
                           n6078);
   U3046 : AO4 port map( A => n4405, B => n7715, C => n2358, D => n7701, Z => 
                           n6079);
   U3047 : AO4 port map( A => n4402, B => n7695, C => n2358, D => n7681, Z => 
                           n6080);
   U3048 : AO4 port map( A => n4403, B => n7675, C => n2358, D => n7661, Z => 
                           n6081);
   U3049 : AO4 port map( A => n4400, B => n7655, C => n2358, D => n7641, Z => 
                           n6082);
   U3050 : AO4 port map( A => n4401, B => n7635, C => n2358, D => n7621, Z => 
                           n6083);
   U3051 : AO4 port map( A => n4398, B => n7615, C => n2357, D => n7601, Z => 
                           n6084);
   U3052 : AO4 port map( A => n4399, B => n7595, C => n2357, D => n7581, Z => 
                           n6085);
   U3053 : AO4 port map( A => n4412, B => n7575, C => n2357, D => n7561, Z => 
                           n6086);
   U3054 : AO4 port map( A => n4413, B => n7555, C => n2357, D => n7541, Z => 
                           n6087);
   U3055 : AO4 port map( A => n4410, B => n7535, C => n2357, D => n7521, Z => 
                           n6088);
   U3056 : AO4 port map( A => n4411, B => n7515, C => n2357, D => n7501, Z => 
                           n6089);
   U3057 : AO4 port map( A => n4408, B => n7495, C => n2357, D => n7481, Z => 
                           n6090);
   U3058 : AO4 port map( A => n4409, B => n7475, C => n2357, D => n7461, Z => 
                           n6091);
   U3059 : AO4 port map( A => n4406, B => n7455, C => n2357, D => n7441, Z => 
                           n6092);
   U3060 : AO4 port map( A => n4407, B => n7435, C => n2357, D => n7421, Z => 
                           n6093);
   U3061 : AO4 port map( A => n4356, B => n7415, C => n2357, D => n7401, Z => 
                           n6094);
   U3062 : AO4 port map( A => n4357, B => n7395, C => n2357, D => n7381, Z => 
                           n6095);
   U3063 : AO4 port map( A => n4354, B => n7375, C => n2357, D => n7361, Z => 
                           n6096);
   U3064 : AO4 port map( A => n4355, B => n7355, C => n2357, D => n7341, Z => 
                           n6097);
   U3065 : AO4 port map( A => n4352, B => n7335, C => n2356, D => n7321, Z => 
                           n6098);
   U3066 : AO4 port map( A => n4353, B => n7315, C => n2356, D => n7301, Z => 
                           n6099);
   U3067 : AO4 port map( A => n4350, B => n7295, C => n2356, D => n7281, Z => 
                           n6100);
   U3068 : AO4 port map( A => n4351, B => n7275, C => n2356, D => n7261, Z => 
                           n6101);
   U3069 : AO4 port map( A => n4364, B => n7255, C => n2356, D => n7241, Z => 
                           n6102);
   U3070 : AO4 port map( A => n4365, B => n7235, C => n2356, D => n7221, Z => 
                           n6103);
   U3071 : AO4 port map( A => n4362, B => n7215, C => n2356, D => n7201, Z => 
                           n6104);
   U3072 : AO4 port map( A => n4363, B => n7195, C => n2356, D => n7181, Z => 
                           n6105);
   U3073 : AO4 port map( A => n4360, B => n7175, C => n2356, D => n7161, Z => 
                           n6106);
   U3074 : AO4 port map( A => n4361, B => n7155, C => n2356, D => n7141, Z => 
                           n6107);
   U3075 : AO4 port map( A => n4358, B => n7135, C => n2356, D => n7121, Z => 
                           n6108);
   U3076 : AO4 port map( A => n4359, B => n7115, C => n2356, D => n7101, Z => 
                           n6109);
   U3077 : AO4 port map( A => n4372, B => n7095, C => n2356, D => n7081, Z => 
                           n6110);
   U3078 : AO4 port map( A => n4373, B => n7075, C => n2356, D => n7061, Z => 
                           n6111);
   U3079 : AO4 port map( A => n4370, B => n7055, C => n2355, D => n7041, Z => 
                           n6112);
   U3080 : AO4 port map( A => n4371, B => n7035, C => n2355, D => n7021, Z => 
                           n6113);
   U3081 : AO4 port map( A => n4368, B => n7015, C => n2355, D => n7001, Z => 
                           n6114);
   U3082 : AO4 port map( A => n4369, B => n6995, C => n2355, D => n6981, Z => 
                           n6115);
   U3083 : AO4 port map( A => n4366, B => n6975, C => n2355, D => n6961, Z => 
                           n6116);
   U3084 : AO4 port map( A => n4367, B => n6955, C => n2355, D => n6941, Z => 
                           n6117);
   U3085 : AO4 port map( A => n4380, B => n6935, C => n2355, D => n6921, Z => 
                           n6118);
   U3086 : AO4 port map( A => n4381, B => n6915, C => n2355, D => n6901, Z => 
                           n6119);
   U3087 : AO4 port map( A => n4378, B => n6895, C => n2355, D => n6881, Z => 
                           n6120);
   U3088 : AO4 port map( A => n4379, B => n6875, C => n2355, D => n6861, Z => 
                           n6121);
   U3089 : AO4 port map( A => n4376, B => n6855, C => n2355, D => n6841, Z => 
                           n6122);
   U3090 : AO4 port map( A => n4377, B => n6835, C => n2355, D => n6821, Z => 
                           n6123);
   U3091 : AO4 port map( A => n4374, B => n6815, C => n2355, D => n6801, Z => 
                           n6124);
   U3092 : AO4 port map( A => n4375, B => n6795, C => n2355, D => n6781, Z => 
                           n6125);
   U3093 : AO4 port map( A => n4460, B => n7896, C => n2310, D => n7877, Z => 
                           n6582);
   U3094 : AO4 port map( A => n4461, B => n7876, C => n2310, D => n7857, Z => 
                           n6583);
   U3095 : AO4 port map( A => n4458, B => n7856, C => n2310, D => n7837, Z => 
                           n6584);
   U3096 : AO4 port map( A => n4459, B => n7836, C => n2310, D => n7817, Z => 
                           n6585);
   U3097 : AO4 port map( A => n4456, B => n7816, C => n2310, D => n7797, Z => 
                           n6586);
   U3098 : AO4 port map( A => n4457, B => n7796, C => n2310, D => n7777, Z => 
                           n6587);
   U3099 : AO4 port map( A => n4454, B => n7776, C => n2310, D => n7757, Z => 
                           n6588);
   U3100 : AO4 port map( A => n4455, B => n7756, C => n2310, D => n7737, Z => 
                           n6589);
   U3101 : AO4 port map( A => n4468, B => n7736, C => n2310, D => n7717, Z => 
                           n6590);
   U3102 : AO4 port map( A => n4469, B => n7716, C => n2310, D => n7697, Z => 
                           n6591);
   U3103 : AO4 port map( A => n4466, B => n7696, C => n2310, D => n7677, Z => 
                           n6592);
   U3104 : AO4 port map( A => n4467, B => n7676, C => n2310, D => n7657, Z => 
                           n6593);
   U3105 : AO4 port map( A => n4464, B => n7656, C => n2310, D => n7637, Z => 
                           n6594);
   U3106 : AO4 port map( A => n4465, B => n7636, C => n2310, D => n7617, Z => 
                           n6595);
   U3107 : AO4 port map( A => n4462, B => n7616, C => n2309, D => n7597, Z => 
                           n6596);
   U3108 : AO4 port map( A => n4463, B => n7596, C => n2309, D => n7577, Z => 
                           n6597);
   U3109 : AO4 port map( A => n4476, B => n7576, C => n2309, D => n7557, Z => 
                           n6598);
   U3110 : AO4 port map( A => n4477, B => n7556, C => n2309, D => n7537, Z => 
                           n6599);
   U3111 : AO4 port map( A => n4474, B => n7536, C => n2309, D => n7517, Z => 
                           n6600);
   U3112 : AO4 port map( A => n4475, B => n7516, C => n2309, D => n7497, Z => 
                           n6601);
   U3113 : AO4 port map( A => n4472, B => n7496, C => n2309, D => n7477, Z => 
                           n6602);
   U3114 : AO4 port map( A => n4473, B => n7476, C => n2309, D => n7457, Z => 
                           n6603);
   U3115 : AO4 port map( A => n4470, B => n7456, C => n2309, D => n7437, Z => 
                           n6604);
   U3116 : AO4 port map( A => n4471, B => n7436, C => n2309, D => n7417, Z => 
                           n6605);
   U3117 : AO4 port map( A => n4420, B => n7416, C => n2309, D => n7397, Z => 
                           n6606);
   U3118 : AO4 port map( A => n4421, B => n7396, C => n2309, D => n7377, Z => 
                           n6607);
   U3119 : AO4 port map( A => n4418, B => n7376, C => n2309, D => n7357, Z => 
                           n6608);
   U3120 : AO4 port map( A => n4419, B => n7356, C => n2309, D => n7337, Z => 
                           n6609);
   U3121 : AO4 port map( A => n4416, B => n7336, C => n2308, D => n7317, Z => 
                           n6610);
   U3122 : AO4 port map( A => n4417, B => n7316, C => n2308, D => n7297, Z => 
                           n6611);
   U3123 : AO4 port map( A => n4414, B => n7296, C => n2308, D => n7277, Z => 
                           n6612);
   U3124 : AO4 port map( A => n4415, B => n7276, C => n2308, D => n7257, Z => 
                           n6613);
   U3125 : AO4 port map( A => n4428, B => n7256, C => n2308, D => n7237, Z => 
                           n6614);
   U3126 : AO4 port map( A => n4429, B => n7236, C => n2308, D => n7217, Z => 
                           n6615);
   U3127 : AO4 port map( A => n4426, B => n7216, C => n2308, D => n7197, Z => 
                           n6616);
   U3128 : AO4 port map( A => n4427, B => n7196, C => n2308, D => n7177, Z => 
                           n6617);
   U3129 : AO4 port map( A => n4424, B => n7176, C => n2308, D => n7157, Z => 
                           n6618);
   U3130 : AO4 port map( A => n4425, B => n7156, C => n2308, D => n7137, Z => 
                           n6619);
   U3131 : AO4 port map( A => n4422, B => n7136, C => n2308, D => n7117, Z => 
                           n6620);
   U3132 : AO4 port map( A => n4423, B => n7116, C => n2308, D => n7097, Z => 
                           n6621);
   U3133 : AO4 port map( A => n4436, B => n7096, C => n2308, D => n7077, Z => 
                           n6622);
   U3134 : AO4 port map( A => n4437, B => n7076, C => n2308, D => n7057, Z => 
                           n6623);
   U3135 : AO4 port map( A => n4434, B => n7056, C => n2307, D => n7037, Z => 
                           n6624);
   U3136 : AO4 port map( A => n4435, B => n7036, C => n2307, D => n7017, Z => 
                           n6625);
   U3137 : AO4 port map( A => n4432, B => n7016, C => n2307, D => n6997, Z => 
                           n6626);
   U3138 : AO4 port map( A => n4433, B => n6996, C => n2307, D => n6977, Z => 
                           n6627);
   U3139 : AO4 port map( A => n4430, B => n6976, C => n2307, D => n6957, Z => 
                           n6628);
   U3140 : AO4 port map( A => n4431, B => n6956, C => n2307, D => n6937, Z => 
                           n6629);
   U3141 : AO4 port map( A => n4444, B => n6936, C => n2307, D => n6917, Z => 
                           n6630);
   U3142 : AO4 port map( A => n4445, B => n6916, C => n2307, D => n6897, Z => 
                           n6631);
   U3143 : AO4 port map( A => n4442, B => n6896, C => n2307, D => n6877, Z => 
                           n6632);
   U3144 : AO4 port map( A => n4443, B => n6876, C => n2307, D => n6857, Z => 
                           n6633);
   U3145 : AO4 port map( A => n4440, B => n6856, C => n2307, D => n6837, Z => 
                           n6634);
   U3146 : AO4 port map( A => n4441, B => n6836, C => n2307, D => n6817, Z => 
                           n6635);
   U3147 : AO4 port map( A => n4438, B => n6816, C => n2307, D => n6797, Z => 
                           n6636);
   U3148 : AO4 port map( A => n4439, B => n6796, C => n2307, D => n6777, Z => 
                           n6637);
   U3149 : AO4 port map( A => n4524, B => n7894, C => n6736, D => n7889, Z => 
                           n5046);
   U3150 : AO4 port map( A => n4525, B => n7874, C => n6736, D => n7869, Z => 
                           n5047);
   U3151 : AO4 port map( A => n4522, B => n7854, C => n6736, D => n7849, Z => 
                           n5048);
   U3152 : AO4 port map( A => n4523, B => n7834, C => n6736, D => n7829, Z => 
                           n5049);
   U3153 : AO4 port map( A => n4520, B => n7814, C => n6736, D => n7809, Z => 
                           n5050);
   U3154 : AO4 port map( A => n4521, B => n7794, C => n6736, D => n7789, Z => 
                           n5051);
   U3155 : AO4 port map( A => n4518, B => n7774, C => n6736, D => n7769, Z => 
                           n5052);
   U3156 : AO4 port map( A => n4519, B => n7754, C => n6736, D => n7749, Z => 
                           n5053);
   U3157 : AO4 port map( A => n4532, B => n7734, C => n6736, D => n7729, Z => 
                           n5054);
   U3158 : AO4 port map( A => n4533, B => n7714, C => n6736, D => n7709, Z => 
                           n5055);
   U3159 : AO4 port map( A => n4530, B => n7694, C => n6736, D => n7689, Z => 
                           n5056);
   U3160 : AO4 port map( A => n4531, B => n7674, C => n6736, D => n7669, Z => 
                           n5057);
   U3161 : AO4 port map( A => n4528, B => n7654, C => n6736, D => n7649, Z => 
                           n5058);
   U3162 : AO4 port map( A => n4529, B => n7634, C => n6736, D => n7629, Z => 
                           n5059);
   U3163 : AO4 port map( A => n4526, B => n7614, C => n6735, D => n7609, Z => 
                           n5060);
   U3164 : AO4 port map( A => n4527, B => n7594, C => n6735, D => n7589, Z => 
                           n5061);
   U3165 : AO4 port map( A => n4540, B => n7574, C => n6735, D => n7569, Z => 
                           n5062);
   U3166 : AO4 port map( A => n4541, B => n7554, C => n6735, D => n7549, Z => 
                           n5063);
   U3167 : AO4 port map( A => n4538, B => n7534, C => n6735, D => n7529, Z => 
                           n5064);
   U3168 : AO4 port map( A => n4539, B => n7514, C => n6735, D => n7509, Z => 
                           n5065);
   U3169 : AO4 port map( A => n4536, B => n7494, C => n6735, D => n7489, Z => 
                           n5066);
   U3170 : AO4 port map( A => n4537, B => n7474, C => n6735, D => n7469, Z => 
                           n5067);
   U3171 : AO4 port map( A => n4534, B => n7454, C => n6735, D => n7449, Z => 
                           n5068);
   U3172 : AO4 port map( A => n4535, B => n7434, C => n6735, D => n7429, Z => 
                           n5069);
   U3173 : AO4 port map( A => n4484, B => n7414, C => n6735, D => n7409, Z => 
                           n5070);
   U3174 : AO4 port map( A => n4485, B => n7394, C => n6735, D => n7389, Z => 
                           n5071);
   U3175 : AO4 port map( A => n4482, B => n7374, C => n6735, D => n7369, Z => 
                           n5072);
   U3176 : AO4 port map( A => n4483, B => n7354, C => n6735, D => n7349, Z => 
                           n5073);
   U3177 : AO4 port map( A => n4480, B => n7334, C => n6734, D => n7329, Z => 
                           n5074);
   U3178 : AO4 port map( A => n4481, B => n7314, C => n6734, D => n7309, Z => 
                           n5075);
   U3179 : AO4 port map( A => n4478, B => n7294, C => n6734, D => n7289, Z => 
                           n5076);
   U3180 : AO4 port map( A => n4479, B => n7274, C => n6734, D => n7269, Z => 
                           n5077);
   U3181 : AO4 port map( A => n4492, B => n7254, C => n6734, D => n7249, Z => 
                           n5078);
   U3182 : AO4 port map( A => n4493, B => n7234, C => n6734, D => n7229, Z => 
                           n5079);
   U3183 : AO4 port map( A => n4490, B => n7214, C => n6734, D => n7209, Z => 
                           n5080);
   U3184 : AO4 port map( A => n4491, B => n7194, C => n6734, D => n7189, Z => 
                           n5081);
   U3185 : AO4 port map( A => n4488, B => n7174, C => n6734, D => n7169, Z => 
                           n5082);
   U3186 : AO4 port map( A => n4489, B => n7154, C => n6734, D => n7149, Z => 
                           n5083);
   U3187 : AO4 port map( A => n4486, B => n7134, C => n6734, D => n7129, Z => 
                           n5084);
   U3188 : AO4 port map( A => n4487, B => n7114, C => n6734, D => n7109, Z => 
                           n5085);
   U3189 : AO4 port map( A => n4500, B => n7094, C => n6734, D => n7089, Z => 
                           n5086);
   U3190 : AO4 port map( A => n4501, B => n7074, C => n6734, D => n7069, Z => 
                           n5087);
   U3191 : AO4 port map( A => n4498, B => n7054, C => n6733, D => n7049, Z => 
                           n5088);
   U3192 : AO4 port map( A => n4499, B => n7034, C => n6733, D => n7029, Z => 
                           n5089);
   U3193 : AO4 port map( A => n4496, B => n7014, C => n6733, D => n7009, Z => 
                           n5090);
   U3194 : AO4 port map( A => n4497, B => n6994, C => n6733, D => n6989, Z => 
                           n5091);
   U3195 : AO4 port map( A => n4494, B => n6974, C => n6733, D => n6969, Z => 
                           n5092);
   U3196 : AO4 port map( A => n4495, B => n6954, C => n6733, D => n6949, Z => 
                           n5093);
   U3197 : AO4 port map( A => n4508, B => n6934, C => n6733, D => n6929, Z => 
                           n5094);
   U3198 : AO4 port map( A => n4509, B => n6914, C => n6733, D => n6909, Z => 
                           n5095);
   U3199 : AO4 port map( A => n4506, B => n6894, C => n6733, D => n6889, Z => 
                           n5096);
   U3200 : AO4 port map( A => n4507, B => n6874, C => n6733, D => n6869, Z => 
                           n5097);
   U3201 : AO4 port map( A => n4504, B => n6854, C => n6733, D => n6849, Z => 
                           n5098);
   U3202 : AO4 port map( A => n4505, B => n6834, C => n6733, D => n6829, Z => 
                           n5099);
   U3203 : AO4 port map( A => n4502, B => n6814, C => n6733, D => n6809, Z => 
                           n5100);
   U3204 : AO4 port map( A => n4503, B => n6794, C => n6733, D => n6789, Z => 
                           n5101);
   U3205 : NR4 port map( A => n347, B => n348, C => n349, D => n350, Z => n346)
                           ;
   U3206 : AO4 port map( A => n2525, B => n8120, C => n2524, D => n8119, Z => 
                           n347);
   U3207 : AO4 port map( A => n2527, B => n8122, C => n2526, D => n8121, Z => 
                           n348);
   U3208 : AO4 port map( A => n2529, B => n8124, C => n2528, D => n8123, Z => 
                           n349);
   U3209 : NR4 port map( A => n359, B => n360, C => n361, D => n362, Z => n345)
                           ;
   U3210 : AO4 port map( A => n2533, B => n8112, C => n2532, D => n8111, Z => 
                           n359);
   U3211 : AO4 port map( A => n2535, B => n8114, C => n2534, D => n8113, Z => 
                           n360);
   U3212 : AO4 port map( A => n2537, B => n8116, C => n2536, D => n8115, Z => 
                           n361);
   U3213 : NR4 port map( A => n371, B => n372, C => n373, D => n374, Z => n344)
                           ;
   U3214 : AO4 port map( A => n2541, B => n8104, C => n2540, D => n8103, Z => 
                           n371);
   U3215 : AO4 port map( A => n2543, B => n8106, C => n2542, D => n8105, Z => 
                           n372);
   U3216 : AO4 port map( A => n2545, B => n8108, C => n2544, D => n8107, Z => 
                           n373);
   U3217 : NR4 port map( A => n383, B => n384, C => n385, D => n386, Z => n343)
                           ;
   U3218 : AO4 port map( A => n2549, B => n8096, C => n2548, D => n8095, Z => 
                           n383);
   U3219 : AO4 port map( A => n2551, B => n8098, C => n2550, D => n8097, Z => 
                           n384);
   U3220 : AO4 port map( A => n2553, B => n8100, C => n2552, D => n8099, Z => 
                           n385);
   U3221 : NR4 port map( A => n399, B => n400, C => n401, D => n402, Z => n398)
                           ;
   U3222 : AO4 port map( A => n2493, B => n8088, C => n2492, D => n8087, Z => 
                           n399);
   U3223 : AO4 port map( A => n2495, B => n8090, C => n2494, D => n8089, Z => 
                           n400);
   U3224 : AO4 port map( A => n2497, B => n8092, C => n2496, D => n8091, Z => 
                           n401);
   U3225 : NR4 port map( A => n411, B => n412, C => n413, D => n414, Z => n397)
                           ;
   U3226 : AO4 port map( A => n2501, B => n8080, C => n2500, D => n8079, Z => 
                           n411);
   U3227 : AO4 port map( A => n2503, B => n8082, C => n2502, D => n8081, Z => 
                           n412);
   U3228 : AO4 port map( A => n2505, B => n8084, C => n2504, D => n8083, Z => 
                           n413);
   U3229 : NR4 port map( A => n423, B => n424, C => n425, D => n426, Z => n396)
                           ;
   U3230 : AO4 port map( A => n2509, B => n8072, C => n2508, D => n8071, Z => 
                           n423);
   U3231 : AO4 port map( A => n2511, B => n8074, C => n2510, D => n8073, Z => 
                           n424);
   U3232 : AO4 port map( A => n2513, B => n8076, C => n2512, D => n8075, Z => 
                           n425);
   U3233 : NR4 port map( A => n435, B => n436, C => n437, D => n438, Z => n395)
                           ;
   U3234 : AO4 port map( A => n2517, B => n8064, C => n2516, D => n8063, Z => 
                           n435);
   U3235 : AO4 port map( A => n2519, B => n8066, C => n2518, D => n8065, Z => 
                           n436);
   U3236 : AO4 port map( A => n2521, B => n8068, C => n2520, D => n8067, Z => 
                           n437);
   U3237 : NR4 port map( A => n455, B => n456, C => n457, D => n458, Z => n454)
                           ;
   U3238 : AO4 port map( A => n2589, B => n8120, C => n2588, D => n8119, Z => 
                           n455);
   U3239 : AO4 port map( A => n2591, B => n8122, C => n2590, D => n8121, Z => 
                           n456);
   U3240 : AO4 port map( A => n2593, B => n8124, C => n2592, D => n8123, Z => 
                           n457);
   U3241 : NR4 port map( A => n459, B => n460, C => n461, D => n462, Z => n453)
                           ;
   U3242 : AO4 port map( A => n2597, B => n8112, C => n2596, D => n8111, Z => 
                           n459);
   U3243 : AO4 port map( A => n2599, B => n8114, C => n2598, D => n8113, Z => 
                           n460);
   U3244 : AO4 port map( A => n2601, B => n8116, C => n2600, D => n8115, Z => 
                           n461);
   U3245 : NR4 port map( A => n463, B => n464, C => n465, D => n466, Z => n452)
                           ;
   U3246 : AO4 port map( A => n2605, B => n8104, C => n2604, D => n8103, Z => 
                           n463);
   U3247 : AO4 port map( A => n2607, B => n8106, C => n2606, D => n8105, Z => 
                           n464);
   U3248 : AO4 port map( A => n2609, B => n8108, C => n2608, D => n8107, Z => 
                           n465);
   U3249 : NR4 port map( A => n467, B => n468, C => n469, D => n470, Z => n451)
                           ;
   U3250 : AO4 port map( A => n2613, B => n8096, C => n2612, D => n8095, Z => 
                           n467);
   U3251 : AO4 port map( A => n2615, B => n8098, C => n2614, D => n8097, Z => 
                           n468);
   U3252 : AO4 port map( A => n2617, B => n8100, C => n2616, D => n8099, Z => 
                           n469);
   U3253 : NR4 port map( A => n475, B => n476, C => n477, D => n478, Z => n474)
                           ;
   U3254 : AO4 port map( A => n2557, B => n8088, C => n2556, D => n8087, Z => 
                           n475);
   U3255 : AO4 port map( A => n2559, B => n8090, C => n2558, D => n8089, Z => 
                           n476);
   U3256 : AO4 port map( A => n2561, B => n8092, C => n2560, D => n8091, Z => 
                           n477);
   U3257 : NR4 port map( A => n479, B => n480, C => n481, D => n482, Z => n473)
                           ;
   U3258 : AO4 port map( A => n2565, B => n8080, C => n2564, D => n8079, Z => 
                           n479);
   U3259 : AO4 port map( A => n2567, B => n8082, C => n2566, D => n8081, Z => 
                           n480);
   U3260 : AO4 port map( A => n2569, B => n8084, C => n2568, D => n8083, Z => 
                           n481);
   U3261 : NR4 port map( A => n483, B => n484, C => n485, D => n486, Z => n472)
                           ;
   U3262 : AO4 port map( A => n2573, B => n8072, C => n2572, D => n8071, Z => 
                           n483);
   U3263 : AO4 port map( A => n2575, B => n8074, C => n2574, D => n8073, Z => 
                           n484);
   U3264 : AO4 port map( A => n2577, B => n8076, C => n2576, D => n8075, Z => 
                           n485);
   U3265 : NR4 port map( A => n487, B => n488, C => n489, D => n490, Z => n471)
                           ;
   U3266 : AO4 port map( A => n2581, B => n8064, C => n2580, D => n8063, Z => 
                           n487);
   U3267 : AO4 port map( A => n2583, B => n8066, C => n2582, D => n8065, Z => 
                           n488);
   U3268 : AO4 port map( A => n2585, B => n8068, C => n2584, D => n8067, Z => 
                           n489);
   U3269 : NR4 port map( A => n499, B => n500, C => n501, D => n502, Z => n498)
                           ;
   U3270 : AO4 port map( A => n2653, B => n8120, C => n2652, D => n8119, Z => 
                           n499);
   U3271 : AO4 port map( A => n2655, B => n8122, C => n2654, D => n8121, Z => 
                           n500);
   U3272 : AO4 port map( A => n2657, B => n8124, C => n2656, D => n8123, Z => 
                           n501);
   U3273 : NR4 port map( A => n503, B => n504, C => n505, D => n506, Z => n497)
                           ;
   U3274 : AO4 port map( A => n2661, B => n8112, C => n2660, D => n8111, Z => 
                           n503);
   U3275 : AO4 port map( A => n2663, B => n8114, C => n2662, D => n8113, Z => 
                           n504);
   U3276 : AO4 port map( A => n2665, B => n8116, C => n2664, D => n8115, Z => 
                           n505);
   U3277 : NR4 port map( A => n507, B => n508, C => n509, D => n510, Z => n496)
                           ;
   U3278 : AO4 port map( A => n2669, B => n8104, C => n2668, D => n8103, Z => 
                           n507);
   U3279 : AO4 port map( A => n2671, B => n8106, C => n2670, D => n8105, Z => 
                           n508);
   U3280 : AO4 port map( A => n2673, B => n8108, C => n2672, D => n8107, Z => 
                           n509);
   U3281 : NR4 port map( A => n511, B => n512, C => n513, D => n514, Z => n495)
                           ;
   U3282 : AO4 port map( A => n2677, B => n8096, C => n2676, D => n8095, Z => 
                           n511);
   U3283 : AO4 port map( A => n2679, B => n8098, C => n2678, D => n8097, Z => 
                           n512);
   U3284 : AO4 port map( A => n2681, B => n8100, C => n2680, D => n8099, Z => 
                           n513);
   U3285 : NR4 port map( A => n519, B => n520, C => n521, D => n522, Z => n518)
                           ;
   U3286 : AO4 port map( A => n2621, B => n8088, C => n2620, D => n8087, Z => 
                           n519);
   U3287 : AO4 port map( A => n2623, B => n8090, C => n2622, D => n8089, Z => 
                           n520);
   U3288 : AO4 port map( A => n2625, B => n8092, C => n2624, D => n8091, Z => 
                           n521);
   U3289 : NR4 port map( A => n523, B => n524, C => n525, D => n526, Z => n517)
                           ;
   U3290 : AO4 port map( A => n2629, B => n8080, C => n2628, D => n8079, Z => 
                           n523);
   U3291 : AO4 port map( A => n2631, B => n8082, C => n2630, D => n8081, Z => 
                           n524);
   U3292 : AO4 port map( A => n2633, B => n8084, C => n2632, D => n8083, Z => 
                           n525);
   U3293 : NR4 port map( A => n527, B => n528, C => n529, D => n530, Z => n516)
                           ;
   U3294 : AO4 port map( A => n2637, B => n8072, C => n2636, D => n8071, Z => 
                           n527);
   U3295 : AO4 port map( A => n2639, B => n8074, C => n2638, D => n8073, Z => 
                           n528);
   U3296 : AO4 port map( A => n2641, B => n8076, C => n2640, D => n8075, Z => 
                           n529);
   U3297 : NR4 port map( A => n531, B => n532, C => n533, D => n534, Z => n515)
                           ;
   U3298 : AO4 port map( A => n2645, B => n8064, C => n2644, D => n8063, Z => 
                           n531);
   U3299 : AO4 port map( A => n2647, B => n8066, C => n2646, D => n8065, Z => 
                           n532);
   U3300 : AO4 port map( A => n2649, B => n8068, C => n2648, D => n8067, Z => 
                           n533);
   U3301 : NR4 port map( A => n543, B => n544, C => n545, D => n546, Z => n542)
                           ;
   U3302 : AO4 port map( A => n2717, B => n8120, C => n2716, D => n8119, Z => 
                           n543);
   U3303 : AO4 port map( A => n2719, B => n8122, C => n2718, D => n8121, Z => 
                           n544);
   U3304 : AO4 port map( A => n2721, B => n8124, C => n2720, D => n8123, Z => 
                           n545);
   U3305 : NR4 port map( A => n547, B => n548, C => n549, D => n550, Z => n541)
                           ;
   U3306 : AO4 port map( A => n2725, B => n8112, C => n2724, D => n8111, Z => 
                           n547);
   U3307 : AO4 port map( A => n2727, B => n8114, C => n2726, D => n8113, Z => 
                           n548);
   U3308 : AO4 port map( A => n2729, B => n8116, C => n2728, D => n8115, Z => 
                           n549);
   U3309 : NR4 port map( A => n551, B => n552, C => n553, D => n554, Z => n540)
                           ;
   U3310 : AO4 port map( A => n2733, B => n8104, C => n2732, D => n8103, Z => 
                           n551);
   U3311 : AO4 port map( A => n2735, B => n8106, C => n2734, D => n8105, Z => 
                           n552);
   U3312 : AO4 port map( A => n2737, B => n8108, C => n2736, D => n8107, Z => 
                           n553);
   U3313 : NR4 port map( A => n555, B => n556, C => n557, D => n558, Z => n539)
                           ;
   U3314 : AO4 port map( A => n2741, B => n8096, C => n2740, D => n8095, Z => 
                           n555);
   U3315 : AO4 port map( A => n2743, B => n8098, C => n2742, D => n8097, Z => 
                           n556);
   U3316 : AO4 port map( A => n2745, B => n8100, C => n2744, D => n8099, Z => 
                           n557);
   U3317 : NR4 port map( A => n563, B => n564, C => n565, D => n566, Z => n562)
                           ;
   U3318 : AO4 port map( A => n2685, B => n8088, C => n2684, D => n8087, Z => 
                           n563);
   U3319 : AO4 port map( A => n2687, B => n8090, C => n2686, D => n8089, Z => 
                           n564);
   U3320 : AO4 port map( A => n2689, B => n8092, C => n2688, D => n8091, Z => 
                           n565);
   U3321 : NR4 port map( A => n567, B => n568, C => n569, D => n570, Z => n561)
                           ;
   U3322 : AO4 port map( A => n2693, B => n8080, C => n2692, D => n8079, Z => 
                           n567);
   U3323 : AO4 port map( A => n2695, B => n8082, C => n2694, D => n8081, Z => 
                           n568);
   U3324 : AO4 port map( A => n2697, B => n8084, C => n2696, D => n8083, Z => 
                           n569);
   U3325 : NR4 port map( A => n571, B => n572, C => n573, D => n574, Z => n560)
                           ;
   U3326 : AO4 port map( A => n2701, B => n8072, C => n2700, D => n8071, Z => 
                           n571);
   U3327 : AO4 port map( A => n2703, B => n8074, C => n2702, D => n8073, Z => 
                           n572);
   U3328 : AO4 port map( A => n2705, B => n8076, C => n2704, D => n8075, Z => 
                           n573);
   U3329 : NR4 port map( A => n575, B => n576, C => n577, D => n578, Z => n559)
                           ;
   U3330 : AO4 port map( A => n2709, B => n8064, C => n2708, D => n8063, Z => 
                           n575);
   U3331 : AO4 port map( A => n2711, B => n8066, C => n2710, D => n8065, Z => 
                           n576);
   U3332 : AO4 port map( A => n2713, B => n8068, C => n2712, D => n8067, Z => 
                           n577);
   U3333 : NR4 port map( A => n587, B => n588, C => n589, D => n590, Z => n586)
                           ;
   U3334 : AO4 port map( A => n2782, B => n8120, C => n2781, D => n8119, Z => 
                           n587);
   U3335 : AO4 port map( A => n2784, B => n8122, C => n2783, D => n8121, Z => 
                           n588);
   U3336 : AO4 port map( A => n2786, B => n8124, C => n2785, D => n8123, Z => 
                           n589);
   U3337 : NR4 port map( A => n591, B => n592, C => n593, D => n594, Z => n585)
                           ;
   U3338 : AO4 port map( A => n2790, B => n8112, C => n2789, D => n8111, Z => 
                           n591);
   U3339 : AO4 port map( A => n2792, B => n8114, C => n2791, D => n8113, Z => 
                           n592);
   U3340 : AO4 port map( A => n2794, B => n8116, C => n2793, D => n8115, Z => 
                           n593);
   U3341 : NR4 port map( A => n595, B => n596, C => n597, D => n598, Z => n584)
                           ;
   U3342 : AO4 port map( A => n2798, B => n8104, C => n2797, D => n8103, Z => 
                           n595);
   U3343 : AO4 port map( A => n2800, B => n8106, C => n2799, D => n8105, Z => 
                           n596);
   U3344 : AO4 port map( A => n2802, B => n8108, C => n2801, D => n8107, Z => 
                           n597);
   U3345 : NR4 port map( A => n599, B => n600, C => n601, D => n602, Z => n583)
                           ;
   U3346 : AO4 port map( A => n2806, B => n8096, C => n2805, D => n8095, Z => 
                           n599);
   U3347 : AO4 port map( A => n2808, B => n8098, C => n2807, D => n8097, Z => 
                           n600);
   U3348 : AO4 port map( A => n2810, B => n8100, C => n2809, D => n8099, Z => 
                           n601);
   U3349 : NR4 port map( A => n607, B => n608, C => n609, D => n610, Z => n606)
                           ;
   U3350 : AO4 port map( A => n2750, B => n8088, C => n2749, D => n8087, Z => 
                           n607);
   U3351 : AO4 port map( A => n2752, B => n8090, C => n2751, D => n8089, Z => 
                           n608);
   U3352 : AO4 port map( A => n2754, B => n8092, C => n2753, D => n8091, Z => 
                           n609);
   U3353 : NR4 port map( A => n611, B => n612, C => n613, D => n614, Z => n605)
                           ;
   U3354 : AO4 port map( A => n2758, B => n8080, C => n2757, D => n8079, Z => 
                           n611);
   U3355 : AO4 port map( A => n2760, B => n8082, C => n2759, D => n8081, Z => 
                           n612);
   U3356 : AO4 port map( A => n2762, B => n8084, C => n2761, D => n8083, Z => 
                           n613);
   U3357 : NR4 port map( A => n615, B => n616, C => n617, D => n618, Z => n604)
                           ;
   U3358 : AO4 port map( A => n2766, B => n8072, C => n2765, D => n8071, Z => 
                           n615);
   U3359 : AO4 port map( A => n2768, B => n8074, C => n2767, D => n8073, Z => 
                           n616);
   U3360 : AO4 port map( A => n2770, B => n8076, C => n2769, D => n8075, Z => 
                           n617);
   U3361 : NR4 port map( A => n619, B => n620, C => n621, D => n622, Z => n603)
                           ;
   U3362 : AO4 port map( A => n2774, B => n8064, C => n2773, D => n8063, Z => 
                           n619);
   U3363 : AO4 port map( A => n2776, B => n8066, C => n2775, D => n8065, Z => 
                           n620);
   U3364 : AO4 port map( A => n2778, B => n8068, C => n2777, D => n8067, Z => 
                           n621);
   U3365 : NR4 port map( A => n631, B => n632, C => n633, D => n634, Z => n630)
                           ;
   U3366 : AO4 port map( A => n2846, B => n8120, C => n2845, D => n8119, Z => 
                           n631);
   U3367 : AO4 port map( A => n2848, B => n8122, C => n2847, D => n8121, Z => 
                           n632);
   U3368 : AO4 port map( A => n2850, B => n8124, C => n2849, D => n8123, Z => 
                           n633);
   U3369 : NR4 port map( A => n635, B => n636, C => n637, D => n638, Z => n629)
                           ;
   U3370 : AO4 port map( A => n2854, B => n8112, C => n2853, D => n8111, Z => 
                           n635);
   U3371 : AO4 port map( A => n2856, B => n8114, C => n2855, D => n8113, Z => 
                           n636);
   U3372 : AO4 port map( A => n2858, B => n8116, C => n2857, D => n8115, Z => 
                           n637);
   U3373 : NR4 port map( A => n639, B => n640, C => n641, D => n642, Z => n628)
                           ;
   U3374 : AO4 port map( A => n2862, B => n8104, C => n2861, D => n8103, Z => 
                           n639);
   U3375 : AO4 port map( A => n2864, B => n8106, C => n2863, D => n8105, Z => 
                           n640);
   U3376 : AO4 port map( A => n2866, B => n8108, C => n2865, D => n8107, Z => 
                           n641);
   U3377 : NR4 port map( A => n643, B => n644, C => n645, D => n646, Z => n627)
                           ;
   U3378 : AO4 port map( A => n2870, B => n8096, C => n2869, D => n8095, Z => 
                           n643);
   U3379 : AO4 port map( A => n2872, B => n8098, C => n2871, D => n8097, Z => 
                           n644);
   U3380 : AO4 port map( A => n2874, B => n8100, C => n2873, D => n8099, Z => 
                           n645);
   U3381 : NR4 port map( A => n651, B => n652, C => n653, D => n654, Z => n650)
                           ;
   U3382 : AO4 port map( A => n2814, B => n8088, C => n2813, D => n8087, Z => 
                           n651);
   U3383 : AO4 port map( A => n2816, B => n8090, C => n2815, D => n8089, Z => 
                           n652);
   U3384 : AO4 port map( A => n2818, B => n8092, C => n2817, D => n8091, Z => 
                           n653);
   U3385 : NR4 port map( A => n655, B => n656, C => n657, D => n658, Z => n649)
                           ;
   U3386 : AO4 port map( A => n2822, B => n8080, C => n2821, D => n8079, Z => 
                           n655);
   U3387 : AO4 port map( A => n2824, B => n8082, C => n2823, D => n8081, Z => 
                           n656);
   U3388 : AO4 port map( A => n2826, B => n8084, C => n2825, D => n8083, Z => 
                           n657);
   U3389 : NR4 port map( A => n659, B => n660, C => n661, D => n662, Z => n648)
                           ;
   U3390 : AO4 port map( A => n2830, B => n8072, C => n2829, D => n8071, Z => 
                           n659);
   U3391 : AO4 port map( A => n2832, B => n8074, C => n2831, D => n8073, Z => 
                           n660);
   U3392 : AO4 port map( A => n2834, B => n8076, C => n2833, D => n8075, Z => 
                           n661);
   U3393 : NR4 port map( A => n663, B => n664, C => n665, D => n666, Z => n647)
                           ;
   U3394 : AO4 port map( A => n2838, B => n8064, C => n2837, D => n8063, Z => 
                           n663);
   U3395 : AO4 port map( A => n2840, B => n8066, C => n2839, D => n8065, Z => 
                           n664);
   U3396 : AO4 port map( A => n2842, B => n8068, C => n2841, D => n8067, Z => 
                           n665);
   U3397 : NR4 port map( A => n675, B => n676, C => n677, D => n678, Z => n674)
                           ;
   U3398 : AO4 port map( A => n2910, B => n8120, C => n2909, D => n8119, Z => 
                           n675);
   U3399 : AO4 port map( A => n2912, B => n8122, C => n2911, D => n8121, Z => 
                           n676);
   U3400 : AO4 port map( A => n2914, B => n8124, C => n2913, D => n8123, Z => 
                           n677);
   U3401 : NR4 port map( A => n679, B => n680, C => n681, D => n682, Z => n673)
                           ;
   U3402 : AO4 port map( A => n2918, B => n8112, C => n2917, D => n8111, Z => 
                           n679);
   U3403 : AO4 port map( A => n2920, B => n8114, C => n2919, D => n8113, Z => 
                           n680);
   U3404 : AO4 port map( A => n2922, B => n8116, C => n2921, D => n8115, Z => 
                           n681);
   U3405 : NR4 port map( A => n683, B => n684, C => n685, D => n686, Z => n672)
                           ;
   U3406 : AO4 port map( A => n2926, B => n8104, C => n2925, D => n8103, Z => 
                           n683);
   U3407 : AO4 port map( A => n2928, B => n8106, C => n2927, D => n8105, Z => 
                           n684);
   U3408 : AO4 port map( A => n2930, B => n8108, C => n2929, D => n8107, Z => 
                           n685);
   U3409 : NR4 port map( A => n687, B => n688, C => n689, D => n690, Z => n671)
                           ;
   U3410 : AO4 port map( A => n2934, B => n8096, C => n2933, D => n8095, Z => 
                           n687);
   U3411 : AO4 port map( A => n2936, B => n8098, C => n2935, D => n8097, Z => 
                           n688);
   U3412 : AO4 port map( A => n2938, B => n8100, C => n2937, D => n8099, Z => 
                           n689);
   U3413 : NR4 port map( A => n695, B => n696, C => n697, D => n698, Z => n694)
                           ;
   U3414 : AO4 port map( A => n2878, B => n8088, C => n2877, D => n8087, Z => 
                           n695);
   U3415 : AO4 port map( A => n2880, B => n8090, C => n2879, D => n8089, Z => 
                           n696);
   U3416 : AO4 port map( A => n2882, B => n8092, C => n2881, D => n8091, Z => 
                           n697);
   U3417 : NR4 port map( A => n699, B => n700, C => n701, D => n702, Z => n693)
                           ;
   U3418 : AO4 port map( A => n2886, B => n8080, C => n2885, D => n8079, Z => 
                           n699);
   U3419 : AO4 port map( A => n2888, B => n8082, C => n2887, D => n8081, Z => 
                           n700);
   U3420 : AO4 port map( A => n2890, B => n8084, C => n2889, D => n8083, Z => 
                           n701);
   U3421 : NR4 port map( A => n703, B => n704, C => n705, D => n706, Z => n692)
                           ;
   U3422 : AO4 port map( A => n2894, B => n8072, C => n2893, D => n8071, Z => 
                           n703);
   U3423 : AO4 port map( A => n2896, B => n8074, C => n2895, D => n8073, Z => 
                           n704);
   U3424 : AO4 port map( A => n2898, B => n8076, C => n2897, D => n8075, Z => 
                           n705);
   U3425 : NR4 port map( A => n707, B => n708, C => n709, D => n710, Z => n691)
                           ;
   U3426 : AO4 port map( A => n2902, B => n8064, C => n2901, D => n8063, Z => 
                           n707);
   U3427 : AO4 port map( A => n2904, B => n8066, C => n2903, D => n8065, Z => 
                           n708);
   U3428 : AO4 port map( A => n2906, B => n8068, C => n2905, D => n8067, Z => 
                           n709);
   U3429 : NR4 port map( A => n718, B => n719, C => n720, D => n721, Z => n717)
                           ;
   U3430 : AO4 port map( A => n2974, B => n8120, C => n2973, D => n8119, Z => 
                           n718);
   U3431 : AO4 port map( A => n2976, B => n8122, C => n2975, D => n8121, Z => 
                           n719);
   U3432 : AO4 port map( A => n2978, B => n8124, C => n2977, D => n8123, Z => 
                           n720);
   U3433 : NR4 port map( A => n722, B => n723, C => n724, D => n725, Z => n716)
                           ;
   U3434 : AO4 port map( A => n2982, B => n8112, C => n2981, D => n8111, Z => 
                           n722);
   U3435 : AO4 port map( A => n2984, B => n8114, C => n2983, D => n8113, Z => 
                           n723);
   U3436 : AO4 port map( A => n2986, B => n8116, C => n2985, D => n8115, Z => 
                           n724);
   U3437 : NR4 port map( A => n726, B => n727, C => n728, D => n729, Z => n715)
                           ;
   U3438 : AO4 port map( A => n2990, B => n8104, C => n2989, D => n8103, Z => 
                           n726);
   U3439 : AO4 port map( A => n2992, B => n8106, C => n2991, D => n8105, Z => 
                           n727);
   U3440 : AO4 port map( A => n2994, B => n8108, C => n2993, D => n8107, Z => 
                           n728);
   U3441 : NR4 port map( A => n730, B => n731, C => n732, D => n733, Z => n714)
                           ;
   U3442 : AO4 port map( A => n2998, B => n8096, C => n2997, D => n8095, Z => 
                           n730);
   U3443 : AO4 port map( A => n3000, B => n8098, C => n2999, D => n8097, Z => 
                           n731);
   U3444 : AO4 port map( A => n3002, B => n8100, C => n3001, D => n8099, Z => 
                           n732);
   U3445 : NR4 port map( A => n738, B => n739, C => n740, D => n741, Z => n737)
                           ;
   U3446 : AO4 port map( A => n2942, B => n8088, C => n2941, D => n8087, Z => 
                           n738);
   U3447 : AO4 port map( A => n2944, B => n8090, C => n2943, D => n8089, Z => 
                           n739);
   U3448 : AO4 port map( A => n2946, B => n8092, C => n2945, D => n8091, Z => 
                           n740);
   U3449 : NR4 port map( A => n742, B => n743, C => n744, D => n745, Z => n736)
                           ;
   U3450 : AO4 port map( A => n2950, B => n8080, C => n2949, D => n8079, Z => 
                           n742);
   U3451 : AO4 port map( A => n2952, B => n8082, C => n2951, D => n8081, Z => 
                           n743);
   U3452 : AO4 port map( A => n2954, B => n8084, C => n2953, D => n8083, Z => 
                           n744);
   U3453 : NR4 port map( A => n746, B => n747, C => n748, D => n749, Z => n735)
                           ;
   U3454 : AO4 port map( A => n2958, B => n8072, C => n2957, D => n8071, Z => 
                           n746);
   U3455 : AO4 port map( A => n2960, B => n8074, C => n2959, D => n8073, Z => 
                           n747);
   U3456 : AO4 port map( A => n2962, B => n8076, C => n2961, D => n8075, Z => 
                           n748);
   U3457 : NR4 port map( A => n750, B => n751, C => n752, D => n753, Z => n734)
                           ;
   U3458 : AO4 port map( A => n2966, B => n8064, C => n2965, D => n8063, Z => 
                           n750);
   U3459 : AO4 port map( A => n2968, B => n8066, C => n2967, D => n8065, Z => 
                           n751);
   U3460 : AO4 port map( A => n2970, B => n8068, C => n2969, D => n8067, Z => 
                           n752);
   U3461 : NR4 port map( A => n762, B => n763, C => n764, D => n765, Z => n761)
                           ;
   U3462 : AO4 port map( A => n3038, B => n8120, C => n3037, D => n8119, Z => 
                           n762);
   U3463 : AO4 port map( A => n3040, B => n8122, C => n3039, D => n8121, Z => 
                           n763);
   U3464 : AO4 port map( A => n3042, B => n8124, C => n3041, D => n8123, Z => 
                           n764);
   U3465 : NR4 port map( A => n766, B => n767, C => n768, D => n769, Z => n760)
                           ;
   U3466 : AO4 port map( A => n3046, B => n8112, C => n3045, D => n8111, Z => 
                           n766);
   U3467 : AO4 port map( A => n3048, B => n8114, C => n3047, D => n8113, Z => 
                           n767);
   U3468 : AO4 port map( A => n3050, B => n8116, C => n3049, D => n8115, Z => 
                           n768);
   U3469 : NR4 port map( A => n770, B => n771, C => n772, D => n773, Z => n759)
                           ;
   U3470 : AO4 port map( A => n3054, B => n8104, C => n3053, D => n8103, Z => 
                           n770);
   U3471 : AO4 port map( A => n3056, B => n8106, C => n3055, D => n8105, Z => 
                           n771);
   U3472 : AO4 port map( A => n3058, B => n8108, C => n3057, D => n8107, Z => 
                           n772);
   U3473 : NR4 port map( A => n774, B => n775, C => n776, D => n777, Z => n758)
                           ;
   U3474 : AO4 port map( A => n3062, B => n8096, C => n3061, D => n8095, Z => 
                           n774);
   U3475 : AO4 port map( A => n3064, B => n8098, C => n3063, D => n8097, Z => 
                           n775);
   U3476 : AO4 port map( A => n3066, B => n8100, C => n3065, D => n8099, Z => 
                           n776);
   U3477 : NR4 port map( A => n782, B => n783, C => n784, D => n785, Z => n781)
                           ;
   U3478 : AO4 port map( A => n3006, B => n8088, C => n3005, D => n8087, Z => 
                           n782);
   U3479 : AO4 port map( A => n3008, B => n8090, C => n3007, D => n8089, Z => 
                           n783);
   U3480 : AO4 port map( A => n3010, B => n8092, C => n3009, D => n8091, Z => 
                           n784);
   U3481 : NR4 port map( A => n786, B => n787, C => n788, D => n789, Z => n780)
                           ;
   U3482 : AO4 port map( A => n3014, B => n8080, C => n3013, D => n8079, Z => 
                           n786);
   U3483 : AO4 port map( A => n3016, B => n8082, C => n3015, D => n8081, Z => 
                           n787);
   U3484 : AO4 port map( A => n3018, B => n8084, C => n3017, D => n8083, Z => 
                           n788);
   U3485 : NR4 port map( A => n790, B => n791, C => n792, D => n793, Z => n779)
                           ;
   U3486 : AO4 port map( A => n3022, B => n8072, C => n3021, D => n8071, Z => 
                           n790);
   U3487 : AO4 port map( A => n3024, B => n8074, C => n3023, D => n8073, Z => 
                           n791);
   U3488 : AO4 port map( A => n3026, B => n8076, C => n3025, D => n8075, Z => 
                           n792);
   U3489 : NR4 port map( A => n794, B => n795, C => n796, D => n797, Z => n778)
                           ;
   U3490 : AO4 port map( A => n3030, B => n8064, C => n3029, D => n8063, Z => 
                           n794);
   U3491 : AO4 port map( A => n3032, B => n8066, C => n3031, D => n8065, Z => 
                           n795);
   U3492 : AO4 port map( A => n3034, B => n8068, C => n3033, D => n8067, Z => 
                           n796);
   U3493 : NR4 port map( A => n806, B => n807, C => n808, D => n809, Z => n805)
                           ;
   U3494 : AO4 port map( A => n3102, B => n8120, C => n3101, D => n8119, Z => 
                           n806);
   U3495 : AO4 port map( A => n3104, B => n8122, C => n3103, D => n8121, Z => 
                           n807);
   U3496 : AO4 port map( A => n3106, B => n8124, C => n3105, D => n8123, Z => 
                           n808);
   U3497 : NR4 port map( A => n810, B => n811, C => n812, D => n813, Z => n804)
                           ;
   U3498 : AO4 port map( A => n3110, B => n8112, C => n3109, D => n8111, Z => 
                           n810);
   U3499 : AO4 port map( A => n3112, B => n8114, C => n3111, D => n8113, Z => 
                           n811);
   U3500 : AO4 port map( A => n3114, B => n8116, C => n3113, D => n8115, Z => 
                           n812);
   U3501 : NR4 port map( A => n814, B => n815, C => n816, D => n817, Z => n803)
                           ;
   U3502 : AO4 port map( A => n3118, B => n8104, C => n3117, D => n8103, Z => 
                           n814);
   U3503 : AO4 port map( A => n3120, B => n8106, C => n3119, D => n8105, Z => 
                           n815);
   U3504 : AO4 port map( A => n3122, B => n8108, C => n3121, D => n8107, Z => 
                           n816);
   U3505 : NR4 port map( A => n818, B => n819, C => n820, D => n821, Z => n802)
                           ;
   U3506 : AO4 port map( A => n3126, B => n8096, C => n3125, D => n8095, Z => 
                           n818);
   U3507 : AO4 port map( A => n3128, B => n8098, C => n3127, D => n8097, Z => 
                           n819);
   U3508 : AO4 port map( A => n3130, B => n8100, C => n3129, D => n8099, Z => 
                           n820);
   U3509 : NR4 port map( A => n826, B => n827, C => n828, D => n829, Z => n825)
                           ;
   U3510 : AO4 port map( A => n3070, B => n8088, C => n3069, D => n8087, Z => 
                           n826);
   U3511 : AO4 port map( A => n3072, B => n8090, C => n3071, D => n8089, Z => 
                           n827);
   U3512 : AO4 port map( A => n3074, B => n8092, C => n3073, D => n8091, Z => 
                           n828);
   U3513 : NR4 port map( A => n830, B => n831, C => n832, D => n833, Z => n824)
                           ;
   U3514 : AO4 port map( A => n3078, B => n8080, C => n3077, D => n8079, Z => 
                           n830);
   U3515 : AO4 port map( A => n3080, B => n8082, C => n3079, D => n8081, Z => 
                           n831);
   U3516 : AO4 port map( A => n3082, B => n8084, C => n3081, D => n8083, Z => 
                           n832);
   U3517 : NR4 port map( A => n834, B => n835, C => n836, D => n837, Z => n823)
                           ;
   U3518 : AO4 port map( A => n3086, B => n8072, C => n3085, D => n8071, Z => 
                           n834);
   U3519 : AO4 port map( A => n3088, B => n8074, C => n3087, D => n8073, Z => 
                           n835);
   U3520 : AO4 port map( A => n3090, B => n8076, C => n3089, D => n8075, Z => 
                           n836);
   U3521 : NR4 port map( A => n838, B => n839, C => n840, D => n841, Z => n822)
                           ;
   U3522 : AO4 port map( A => n3094, B => n8064, C => n3093, D => n8063, Z => 
                           n838);
   U3523 : AO4 port map( A => n3096, B => n8066, C => n3095, D => n8065, Z => 
                           n839);
   U3524 : AO4 port map( A => n3098, B => n8068, C => n3097, D => n8067, Z => 
                           n840);
   U3525 : NR4 port map( A => n850, B => n851, C => n852, D => n853, Z => n849)
                           ;
   U3526 : AO4 port map( A => n3166, B => n8120, C => n3165, D => n8119, Z => 
                           n850);
   U3527 : AO4 port map( A => n3168, B => n8122, C => n3167, D => n8121, Z => 
                           n851);
   U3528 : AO4 port map( A => n3170, B => n8124, C => n3169, D => n8123, Z => 
                           n852);
   U3529 : NR4 port map( A => n854, B => n855, C => n856, D => n857, Z => n848)
                           ;
   U3530 : AO4 port map( A => n3174, B => n8112, C => n3173, D => n8111, Z => 
                           n854);
   U3531 : AO4 port map( A => n3176, B => n8114, C => n3175, D => n8113, Z => 
                           n855);
   U3532 : AO4 port map( A => n3178, B => n8116, C => n3177, D => n8115, Z => 
                           n856);
   U3533 : NR4 port map( A => n858, B => n859, C => n860, D => n861, Z => n847)
                           ;
   U3534 : AO4 port map( A => n3182, B => n8104, C => n3181, D => n8103, Z => 
                           n858);
   U3535 : AO4 port map( A => n3184, B => n8106, C => n3183, D => n8105, Z => 
                           n859);
   U3536 : AO4 port map( A => n3186, B => n8108, C => n3185, D => n8107, Z => 
                           n860);
   U3537 : NR4 port map( A => n862, B => n863, C => n864, D => n865, Z => n846)
                           ;
   U3538 : AO4 port map( A => n3190, B => n8096, C => n3189, D => n8095, Z => 
                           n862);
   U3539 : AO4 port map( A => n3192, B => n8098, C => n3191, D => n8097, Z => 
                           n863);
   U3540 : AO4 port map( A => n3194, B => n8100, C => n3193, D => n8099, Z => 
                           n864);
   U3541 : NR4 port map( A => n870, B => n871, C => n872, D => n873, Z => n869)
                           ;
   U3542 : AO4 port map( A => n3134, B => n8088, C => n3133, D => n8087, Z => 
                           n870);
   U3543 : AO4 port map( A => n3136, B => n8090, C => n3135, D => n8089, Z => 
                           n871);
   U3544 : AO4 port map( A => n3138, B => n8092, C => n3137, D => n8091, Z => 
                           n872);
   U3545 : NR4 port map( A => n874, B => n875, C => n876, D => n877, Z => n868)
                           ;
   U3546 : AO4 port map( A => n3142, B => n8080, C => n3141, D => n8079, Z => 
                           n874);
   U3547 : AO4 port map( A => n3144, B => n8082, C => n3143, D => n8081, Z => 
                           n875);
   U3548 : AO4 port map( A => n3146, B => n8084, C => n3145, D => n8083, Z => 
                           n876);
   U3549 : NR4 port map( A => n878, B => n879, C => n880, D => n881, Z => n867)
                           ;
   U3550 : AO4 port map( A => n3150, B => n8072, C => n3149, D => n8071, Z => 
                           n878);
   U3551 : AO4 port map( A => n3152, B => n8074, C => n3151, D => n8073, Z => 
                           n879);
   U3552 : AO4 port map( A => n3154, B => n8076, C => n3153, D => n8075, Z => 
                           n880);
   U3553 : NR4 port map( A => n882, B => n883, C => n884, D => n885, Z => n866)
                           ;
   U3554 : AO4 port map( A => n3158, B => n8064, C => n3157, D => n8063, Z => 
                           n882);
   U3555 : AO4 port map( A => n3160, B => n8066, C => n3159, D => n8065, Z => 
                           n883);
   U3556 : AO4 port map( A => n3162, B => n8068, C => n3161, D => n8067, Z => 
                           n884);
   U3557 : NR4 port map( A => n893, B => n894, C => n895, D => n896, Z => n892)
                           ;
   U3558 : AO4 port map( A => n3230, B => n8120, C => n3229, D => n8119, Z => 
                           n893);
   U3559 : AO4 port map( A => n3232, B => n8122, C => n3231, D => n8121, Z => 
                           n894);
   U3560 : AO4 port map( A => n3234, B => n8124, C => n3233, D => n8123, Z => 
                           n895);
   U3561 : NR4 port map( A => n897, B => n898, C => n899, D => n900, Z => n891)
                           ;
   U3562 : AO4 port map( A => n3238, B => n8112, C => n3237, D => n8111, Z => 
                           n897);
   U3563 : AO4 port map( A => n3240, B => n8114, C => n3239, D => n8113, Z => 
                           n898);
   U3564 : AO4 port map( A => n3242, B => n8116, C => n3241, D => n8115, Z => 
                           n899);
   U3565 : NR4 port map( A => n901, B => n902, C => n903, D => n904, Z => n890)
                           ;
   U3566 : AO4 port map( A => n3246, B => n8104, C => n3245, D => n8103, Z => 
                           n901);
   U3567 : AO4 port map( A => n3248, B => n8106, C => n3247, D => n8105, Z => 
                           n902);
   U3568 : AO4 port map( A => n3250, B => n8108, C => n3249, D => n8107, Z => 
                           n903);
   U3569 : NR4 port map( A => n905, B => n906, C => n907, D => n908, Z => n889)
                           ;
   U3570 : AO4 port map( A => n3254, B => n8096, C => n3253, D => n8095, Z => 
                           n905);
   U3571 : AO4 port map( A => n3256, B => n8098, C => n3255, D => n8097, Z => 
                           n906);
   U3572 : AO4 port map( A => n3258, B => n8100, C => n3257, D => n8099, Z => 
                           n907);
   U3573 : NR4 port map( A => n913, B => n914, C => n915, D => n916, Z => n912)
                           ;
   U3574 : AO4 port map( A => n3198, B => n8088, C => n3197, D => n8087, Z => 
                           n913);
   U3575 : AO4 port map( A => n3200, B => n8090, C => n3199, D => n8089, Z => 
                           n914);
   U3576 : AO4 port map( A => n3202, B => n8092, C => n3201, D => n8091, Z => 
                           n915);
   U3577 : NR4 port map( A => n917, B => n918, C => n919, D => n920, Z => n911)
                           ;
   U3578 : AO4 port map( A => n3206, B => n8080, C => n3205, D => n8079, Z => 
                           n917);
   U3579 : AO4 port map( A => n3208, B => n8082, C => n3207, D => n8081, Z => 
                           n918);
   U3580 : AO4 port map( A => n3210, B => n8084, C => n3209, D => n8083, Z => 
                           n919);
   U3581 : NR4 port map( A => n921, B => n922, C => n923, D => n924, Z => n910)
                           ;
   U3582 : AO4 port map( A => n3214, B => n8072, C => n3213, D => n8071, Z => 
                           n921);
   U3583 : AO4 port map( A => n3216, B => n8074, C => n3215, D => n8073, Z => 
                           n922);
   U3584 : AO4 port map( A => n3218, B => n8076, C => n3217, D => n8075, Z => 
                           n923);
   U3585 : NR4 port map( A => n925, B => n926, C => n927, D => n928, Z => n909)
                           ;
   U3586 : AO4 port map( A => n3222, B => n8064, C => n3221, D => n8063, Z => 
                           n925);
   U3587 : AO4 port map( A => n3224, B => n8066, C => n3223, D => n8065, Z => 
                           n926);
   U3588 : AO4 port map( A => n3226, B => n8068, C => n3225, D => n8067, Z => 
                           n927);
   U3589 : NR4 port map( A => n937, B => n938, C => n939, D => n940, Z => n936)
                           ;
   U3590 : AO4 port map( A => n3294, B => n8120, C => n3293, D => n8119, Z => 
                           n937);
   U3591 : AO4 port map( A => n3296, B => n8122, C => n3295, D => n8121, Z => 
                           n938);
   U3592 : AO4 port map( A => n3298, B => n8124, C => n3297, D => n8123, Z => 
                           n939);
   U3593 : NR4 port map( A => n941, B => n942, C => n943, D => n944, Z => n935)
                           ;
   U3594 : AO4 port map( A => n3302, B => n8112, C => n3301, D => n8111, Z => 
                           n941);
   U3595 : AO4 port map( A => n3304, B => n8114, C => n3303, D => n8113, Z => 
                           n942);
   U3596 : AO4 port map( A => n3306, B => n8116, C => n3305, D => n8115, Z => 
                           n943);
   U3597 : NR4 port map( A => n945, B => n946, C => n947, D => n948, Z => n934)
                           ;
   U3598 : AO4 port map( A => n3310, B => n8104, C => n3309, D => n8103, Z => 
                           n945);
   U3599 : AO4 port map( A => n3312, B => n8106, C => n3311, D => n8105, Z => 
                           n946);
   U3600 : AO4 port map( A => n3314, B => n8108, C => n3313, D => n8107, Z => 
                           n947);
   U3601 : NR4 port map( A => n949, B => n950, C => n951, D => n952, Z => n933)
                           ;
   U3602 : AO4 port map( A => n3318, B => n8096, C => n3317, D => n8095, Z => 
                           n949);
   U3603 : AO4 port map( A => n3320, B => n8098, C => n3319, D => n8097, Z => 
                           n950);
   U3604 : AO4 port map( A => n3322, B => n8100, C => n3321, D => n8099, Z => 
                           n951);
   U3605 : NR4 port map( A => n957, B => n958, C => n959, D => n960, Z => n956)
                           ;
   U3606 : AO4 port map( A => n3262, B => n8088, C => n3261, D => n8087, Z => 
                           n957);
   U3607 : AO4 port map( A => n3264, B => n8090, C => n3263, D => n8089, Z => 
                           n958);
   U3608 : AO4 port map( A => n3266, B => n8092, C => n3265, D => n8091, Z => 
                           n959);
   U3609 : NR4 port map( A => n961, B => n962, C => n963, D => n964, Z => n955)
                           ;
   U3610 : AO4 port map( A => n3270, B => n8080, C => n3269, D => n8079, Z => 
                           n961);
   U3611 : AO4 port map( A => n3272, B => n8082, C => n3271, D => n8081, Z => 
                           n962);
   U3612 : AO4 port map( A => n3274, B => n8084, C => n3273, D => n8083, Z => 
                           n963);
   U3613 : NR4 port map( A => n965, B => n966, C => n967, D => n968, Z => n954)
                           ;
   U3614 : AO4 port map( A => n3278, B => n8072, C => n3277, D => n8071, Z => 
                           n965);
   U3615 : AO4 port map( A => n3280, B => n8074, C => n3279, D => n8073, Z => 
                           n966);
   U3616 : AO4 port map( A => n3282, B => n8076, C => n3281, D => n8075, Z => 
                           n967);
   U3617 : NR4 port map( A => n969, B => n970, C => n971, D => n972, Z => n953)
                           ;
   U3618 : AO4 port map( A => n3286, B => n8064, C => n3285, D => n8063, Z => 
                           n969);
   U3619 : AO4 port map( A => n3288, B => n8066, C => n3287, D => n8065, Z => 
                           n970);
   U3620 : AO4 port map( A => n3290, B => n8068, C => n3289, D => n8067, Z => 
                           n971);
   U3621 : NR4 port map( A => n981, B => n982, C => n983, D => n984, Z => n980)
                           ;
   U3622 : AO4 port map( A => n3358, B => n8120, C => n3357, D => n8119, Z => 
                           n981);
   U3623 : AO4 port map( A => n3360, B => n8122, C => n3359, D => n8121, Z => 
                           n982);
   U3624 : AO4 port map( A => n3362, B => n8124, C => n3361, D => n8123, Z => 
                           n983);
   U3625 : NR4 port map( A => n985, B => n986, C => n987, D => n988, Z => n979)
                           ;
   U3626 : AO4 port map( A => n3366, B => n8112, C => n3365, D => n8111, Z => 
                           n985);
   U3627 : AO4 port map( A => n3368, B => n8114, C => n3367, D => n8113, Z => 
                           n986);
   U3628 : AO4 port map( A => n3370, B => n8116, C => n3369, D => n8115, Z => 
                           n987);
   U3629 : NR4 port map( A => n989, B => n990, C => n991, D => n992, Z => n978)
                           ;
   U3630 : AO4 port map( A => n3374, B => n8104, C => n3373, D => n8103, Z => 
                           n989);
   U3631 : AO4 port map( A => n3376, B => n8106, C => n3375, D => n8105, Z => 
                           n990);
   U3632 : AO4 port map( A => n3378, B => n8108, C => n3377, D => n8107, Z => 
                           n991);
   U3633 : NR4 port map( A => n993, B => n994, C => n995, D => n996, Z => n977)
                           ;
   U3634 : AO4 port map( A => n3382, B => n8096, C => n3381, D => n8095, Z => 
                           n993);
   U3635 : AO4 port map( A => n3384, B => n8098, C => n3383, D => n8097, Z => 
                           n994);
   U3636 : AO4 port map( A => n3386, B => n8100, C => n3385, D => n8099, Z => 
                           n995);
   U3637 : NR4 port map( A => n1001, B => n1002, C => n1003, D => n1004, Z => 
                           n1000);
   U3638 : AO4 port map( A => n3326, B => n8088, C => n3325, D => n8087, Z => 
                           n1001);
   U3639 : AO4 port map( A => n3328, B => n8090, C => n3327, D => n8089, Z => 
                           n1002);
   U3640 : AO4 port map( A => n3330, B => n8092, C => n3329, D => n8091, Z => 
                           n1003);
   U3641 : NR4 port map( A => n1005, B => n1006, C => n1007, D => n1008, Z => 
                           n999);
   U3642 : AO4 port map( A => n3334, B => n8080, C => n3333, D => n8079, Z => 
                           n1005);
   U3643 : AO4 port map( A => n3336, B => n8082, C => n3335, D => n8081, Z => 
                           n1006);
   U3644 : AO4 port map( A => n3338, B => n8084, C => n3337, D => n8083, Z => 
                           n1007);
   U3645 : NR4 port map( A => n1009, B => n1010, C => n1011, D => n1012, Z => 
                           n998);
   U3646 : AO4 port map( A => n3342, B => n8072, C => n3341, D => n8071, Z => 
                           n1009);
   U3647 : AO4 port map( A => n3344, B => n8074, C => n3343, D => n8073, Z => 
                           n1010);
   U3648 : AO4 port map( A => n3346, B => n8076, C => n3345, D => n8075, Z => 
                           n1011);
   U3649 : NR4 port map( A => n1013, B => n1014, C => n1015, D => n1016, Z => 
                           n997);
   U3650 : AO4 port map( A => n3350, B => n8064, C => n3349, D => n8063, Z => 
                           n1013);
   U3651 : AO4 port map( A => n3352, B => n8066, C => n3351, D => n8065, Z => 
                           n1014);
   U3652 : AO4 port map( A => n3354, B => n8068, C => n3353, D => n8067, Z => 
                           n1015);
   U3653 : NR4 port map( A => n1025, B => n1026, C => n1027, D => n1028, Z => 
                           n1024);
   U3654 : AO4 port map( A => n3422, B => n8120, C => n3421, D => n8119, Z => 
                           n1025);
   U3655 : AO4 port map( A => n3424, B => n8122, C => n3423, D => n8121, Z => 
                           n1026);
   U3656 : AO4 port map( A => n3426, B => n8124, C => n3425, D => n8123, Z => 
                           n1027);
   U3657 : NR4 port map( A => n1029, B => n1030, C => n1031, D => n1032, Z => 
                           n1023);
   U3658 : AO4 port map( A => n3430, B => n8112, C => n3429, D => n8111, Z => 
                           n1029);
   U3659 : AO4 port map( A => n3432, B => n8114, C => n3431, D => n8113, Z => 
                           n1030);
   U3660 : AO4 port map( A => n3434, B => n8116, C => n3433, D => n8115, Z => 
                           n1031);
   U3661 : NR4 port map( A => n1033, B => n1034, C => n1035, D => n1036, Z => 
                           n1022);
   U3662 : AO4 port map( A => n3438, B => n8104, C => n3437, D => n8103, Z => 
                           n1033);
   U3663 : AO4 port map( A => n3440, B => n8106, C => n3439, D => n8105, Z => 
                           n1034);
   U3664 : AO4 port map( A => n3442, B => n8108, C => n3441, D => n8107, Z => 
                           n1035);
   U3665 : NR4 port map( A => n1037, B => n1038, C => n1039, D => n1040, Z => 
                           n1021);
   U3666 : AO4 port map( A => n3446, B => n8096, C => n3445, D => n8095, Z => 
                           n1037);
   U3667 : AO4 port map( A => n3448, B => n8098, C => n3447, D => n8097, Z => 
                           n1038);
   U3668 : AO4 port map( A => n3450, B => n8100, C => n3449, D => n8099, Z => 
                           n1039);
   U3669 : NR4 port map( A => n1045, B => n1046, C => n1047, D => n1048, Z => 
                           n1044);
   U3670 : AO4 port map( A => n3390, B => n8088, C => n3389, D => n8087, Z => 
                           n1045);
   U3671 : AO4 port map( A => n3392, B => n8090, C => n3391, D => n8089, Z => 
                           n1046);
   U3672 : AO4 port map( A => n3394, B => n8092, C => n3393, D => n8091, Z => 
                           n1047);
   U3673 : NR4 port map( A => n1049, B => n1050, C => n1051, D => n1052, Z => 
                           n1043);
   U3674 : AO4 port map( A => n3398, B => n8080, C => n3397, D => n8079, Z => 
                           n1049);
   U3675 : AO4 port map( A => n3400, B => n8082, C => n3399, D => n8081, Z => 
                           n1050);
   U3676 : AO4 port map( A => n3402, B => n8084, C => n3401, D => n8083, Z => 
                           n1051);
   U3677 : NR4 port map( A => n1053, B => n1054, C => n1055, D => n1056, Z => 
                           n1042);
   U3678 : AO4 port map( A => n3406, B => n8072, C => n3405, D => n8071, Z => 
                           n1053);
   U3679 : AO4 port map( A => n3408, B => n8074, C => n3407, D => n8073, Z => 
                           n1054);
   U3680 : AO4 port map( A => n3410, B => n8076, C => n3409, D => n8075, Z => 
                           n1055);
   U3681 : NR4 port map( A => n1057, B => n1058, C => n1059, D => n1060, Z => 
                           n1041);
   U3682 : AO4 port map( A => n3414, B => n8064, C => n3413, D => n8063, Z => 
                           n1057);
   U3683 : AO4 port map( A => n3416, B => n8066, C => n3415, D => n8065, Z => 
                           n1058);
   U3684 : AO4 port map( A => n3418, B => n8068, C => n3417, D => n8067, Z => 
                           n1059);
   U3685 : NR4 port map( A => n1068, B => n1069, C => n1070, D => n1071, Z => 
                           n1067);
   U3686 : AO4 port map( A => n3486, B => n8120, C => n3485, D => n8119, Z => 
                           n1068);
   U3687 : AO4 port map( A => n3488, B => n8122, C => n3487, D => n8121, Z => 
                           n1069);
   U3688 : AO4 port map( A => n3490, B => n8124, C => n3489, D => n8123, Z => 
                           n1070);
   U3689 : NR4 port map( A => n1072, B => n1073, C => n1074, D => n1075, Z => 
                           n1066);
   U3690 : AO4 port map( A => n3494, B => n8112, C => n3493, D => n8111, Z => 
                           n1072);
   U3691 : AO4 port map( A => n3496, B => n8114, C => n3495, D => n8113, Z => 
                           n1073);
   U3692 : AO4 port map( A => n3498, B => n8116, C => n3497, D => n8115, Z => 
                           n1074);
   U3693 : NR4 port map( A => n1076, B => n1077, C => n1078, D => n1079, Z => 
                           n1065);
   U3694 : AO4 port map( A => n3502, B => n8104, C => n3501, D => n8103, Z => 
                           n1076);
   U3695 : AO4 port map( A => n3504, B => n8106, C => n3503, D => n8105, Z => 
                           n1077);
   U3696 : AO4 port map( A => n3506, B => n8108, C => n3505, D => n8107, Z => 
                           n1078);
   U3697 : NR4 port map( A => n1080, B => n1081, C => n1082, D => n1083, Z => 
                           n1064);
   U3698 : AO4 port map( A => n3510, B => n8096, C => n3509, D => n8095, Z => 
                           n1080);
   U3699 : AO4 port map( A => n3512, B => n8098, C => n3511, D => n8097, Z => 
                           n1081);
   U3700 : AO4 port map( A => n3514, B => n8100, C => n3513, D => n8099, Z => 
                           n1082);
   U3701 : NR4 port map( A => n1088, B => n1089, C => n1090, D => n1091, Z => 
                           n1087);
   U3702 : AO4 port map( A => n3454, B => n8088, C => n3453, D => n8087, Z => 
                           n1088);
   U3703 : AO4 port map( A => n3456, B => n8090, C => n3455, D => n8089, Z => 
                           n1089);
   U3704 : AO4 port map( A => n3458, B => n8092, C => n3457, D => n8091, Z => 
                           n1090);
   U3705 : NR4 port map( A => n1092, B => n1093, C => n1094, D => n1095, Z => 
                           n1086);
   U3706 : AO4 port map( A => n3462, B => n8080, C => n3461, D => n8079, Z => 
                           n1092);
   U3707 : AO4 port map( A => n3464, B => n8082, C => n3463, D => n8081, Z => 
                           n1093);
   U3708 : AO4 port map( A => n3466, B => n8084, C => n3465, D => n8083, Z => 
                           n1094);
   U3709 : NR4 port map( A => n1096, B => n1097, C => n1098, D => n1099, Z => 
                           n1085);
   U3710 : AO4 port map( A => n3470, B => n8072, C => n3469, D => n8071, Z => 
                           n1096);
   U3711 : AO4 port map( A => n3472, B => n8074, C => n3471, D => n8073, Z => 
                           n1097);
   U3712 : AO4 port map( A => n3474, B => n8076, C => n3473, D => n8075, Z => 
                           n1098);
   U3713 : NR4 port map( A => n1100, B => n1101, C => n1102, D => n1103, Z => 
                           n1084);
   U3714 : AO4 port map( A => n3478, B => n8064, C => n3477, D => n8063, Z => 
                           n1100);
   U3715 : AO4 port map( A => n3480, B => n8066, C => n3479, D => n8065, Z => 
                           n1101);
   U3716 : AO4 port map( A => n3482, B => n8068, C => n3481, D => n8067, Z => 
                           n1102);
   U3717 : NR4 port map( A => n1112, B => n1113, C => n1114, D => n1115, Z => 
                           n1111);
   U3718 : AO4 port map( A => n3550, B => n8120, C => n3549, D => n8119, Z => 
                           n1112);
   U3719 : AO4 port map( A => n3552, B => n8122, C => n3551, D => n8121, Z => 
                           n1113);
   U3720 : AO4 port map( A => n3554, B => n8124, C => n3553, D => n8123, Z => 
                           n1114);
   U3721 : NR4 port map( A => n1116, B => n1117, C => n1118, D => n1119, Z => 
                           n1110);
   U3722 : AO4 port map( A => n3558, B => n8112, C => n3557, D => n8111, Z => 
                           n1116);
   U3723 : AO4 port map( A => n3560, B => n8114, C => n3559, D => n8113, Z => 
                           n1117);
   U3724 : AO4 port map( A => n3562, B => n8116, C => n3561, D => n8115, Z => 
                           n1118);
   U3725 : NR4 port map( A => n1120, B => n1121, C => n1122, D => n1123, Z => 
                           n1109);
   U3726 : AO4 port map( A => n3566, B => n8104, C => n3565, D => n8103, Z => 
                           n1120);
   U3727 : AO4 port map( A => n3568, B => n8106, C => n3567, D => n8105, Z => 
                           n1121);
   U3728 : AO4 port map( A => n3570, B => n8108, C => n3569, D => n8107, Z => 
                           n1122);
   U3729 : NR4 port map( A => n1124, B => n1125, C => n1126, D => n1127, Z => 
                           n1108);
   U3730 : AO4 port map( A => n3574, B => n8096, C => n3573, D => n8095, Z => 
                           n1124);
   U3731 : AO4 port map( A => n3576, B => n8098, C => n3575, D => n8097, Z => 
                           n1125);
   U3732 : AO4 port map( A => n3578, B => n8100, C => n3577, D => n8099, Z => 
                           n1126);
   U3733 : NR4 port map( A => n1132, B => n1133, C => n1134, D => n1135, Z => 
                           n1131);
   U3734 : AO4 port map( A => n3518, B => n8088, C => n3517, D => n8087, Z => 
                           n1132);
   U3735 : AO4 port map( A => n3520, B => n8090, C => n3519, D => n8089, Z => 
                           n1133);
   U3736 : AO4 port map( A => n3522, B => n8092, C => n3521, D => n8091, Z => 
                           n1134);
   U3737 : NR4 port map( A => n1136, B => n1137, C => n1138, D => n1139, Z => 
                           n1130);
   U3738 : AO4 port map( A => n3526, B => n8080, C => n3525, D => n8079, Z => 
                           n1136);
   U3739 : AO4 port map( A => n3528, B => n8082, C => n3527, D => n8081, Z => 
                           n1137);
   U3740 : AO4 port map( A => n3530, B => n8084, C => n3529, D => n8083, Z => 
                           n1138);
   U3741 : NR4 port map( A => n1140, B => n1141, C => n1142, D => n1143, Z => 
                           n1129);
   U3742 : AO4 port map( A => n3534, B => n8072, C => n3533, D => n8071, Z => 
                           n1140);
   U3743 : AO4 port map( A => n3536, B => n8074, C => n3535, D => n8073, Z => 
                           n1141);
   U3744 : AO4 port map( A => n3538, B => n8076, C => n3537, D => n8075, Z => 
                           n1142);
   U3745 : NR4 port map( A => n1144, B => n1145, C => n1146, D => n1147, Z => 
                           n1128);
   U3746 : AO4 port map( A => n3542, B => n8064, C => n3541, D => n8063, Z => 
                           n1144);
   U3747 : AO4 port map( A => n3544, B => n8066, C => n3543, D => n8065, Z => 
                           n1145);
   U3748 : AO4 port map( A => n3546, B => n8068, C => n3545, D => n8067, Z => 
                           n1146);
   U3749 : NR4 port map( A => n1156, B => n1157, C => n1158, D => n1159, Z => 
                           n1155);
   U3750 : AO4 port map( A => n3614, B => n8120, C => n3613, D => n8119, Z => 
                           n1156);
   U3751 : AO4 port map( A => n3616, B => n8122, C => n3615, D => n8121, Z => 
                           n1157);
   U3752 : AO4 port map( A => n3618, B => n8124, C => n3617, D => n8123, Z => 
                           n1158);
   U3753 : NR4 port map( A => n1160, B => n1161, C => n1162, D => n1163, Z => 
                           n1154);
   U3754 : AO4 port map( A => n3622, B => n8112, C => n3621, D => n8111, Z => 
                           n1160);
   U3755 : AO4 port map( A => n3624, B => n8114, C => n3623, D => n8113, Z => 
                           n1161);
   U3756 : AO4 port map( A => n3626, B => n8116, C => n3625, D => n8115, Z => 
                           n1162);
   U3757 : NR4 port map( A => n1164, B => n1165, C => n1166, D => n1167, Z => 
                           n1153);
   U3758 : AO4 port map( A => n3630, B => n8104, C => n3629, D => n8103, Z => 
                           n1164);
   U3759 : AO4 port map( A => n3632, B => n8106, C => n3631, D => n8105, Z => 
                           n1165);
   U3760 : AO4 port map( A => n3634, B => n8108, C => n3633, D => n8107, Z => 
                           n1166);
   U3761 : NR4 port map( A => n1168, B => n1169, C => n1170, D => n1171, Z => 
                           n1152);
   U3762 : AO4 port map( A => n3638, B => n8096, C => n3637, D => n8095, Z => 
                           n1168);
   U3763 : AO4 port map( A => n3640, B => n8098, C => n3639, D => n8097, Z => 
                           n1169);
   U3764 : AO4 port map( A => n3642, B => n8100, C => n3641, D => n8099, Z => 
                           n1170);
   U3765 : NR4 port map( A => n1176, B => n1177, C => n1178, D => n1179, Z => 
                           n1175);
   U3766 : AO4 port map( A => n3582, B => n8088, C => n3581, D => n8087, Z => 
                           n1176);
   U3767 : AO4 port map( A => n3584, B => n8090, C => n3583, D => n8089, Z => 
                           n1177);
   U3768 : AO4 port map( A => n3586, B => n8092, C => n3585, D => n8091, Z => 
                           n1178);
   U3769 : NR4 port map( A => n1180, B => n1181, C => n1182, D => n1183, Z => 
                           n1174);
   U3770 : AO4 port map( A => n3590, B => n8080, C => n3589, D => n8079, Z => 
                           n1180);
   U3771 : AO4 port map( A => n3592, B => n8082, C => n3591, D => n8081, Z => 
                           n1181);
   U3772 : AO4 port map( A => n3594, B => n8084, C => n3593, D => n8083, Z => 
                           n1182);
   U3773 : NR4 port map( A => n1184, B => n1185, C => n1186, D => n1187, Z => 
                           n1173);
   U3774 : AO4 port map( A => n3598, B => n8072, C => n3597, D => n8071, Z => 
                           n1184);
   U3775 : AO4 port map( A => n3600, B => n8074, C => n3599, D => n8073, Z => 
                           n1185);
   U3776 : AO4 port map( A => n3602, B => n8076, C => n3601, D => n8075, Z => 
                           n1186);
   U3777 : NR4 port map( A => n1188, B => n1189, C => n1190, D => n1191, Z => 
                           n1172);
   U3778 : AO4 port map( A => n3606, B => n8064, C => n3605, D => n8063, Z => 
                           n1188);
   U3779 : AO4 port map( A => n3608, B => n8066, C => n3607, D => n8065, Z => 
                           n1189);
   U3780 : AO4 port map( A => n3610, B => n8068, C => n3609, D => n8067, Z => 
                           n1190);
   U3781 : NR4 port map( A => n1200, B => n1201, C => n1202, D => n1203, Z => 
                           n1199);
   U3782 : AO4 port map( A => n3678, B => n8120, C => n3677, D => n8119, Z => 
                           n1200);
   U3783 : AO4 port map( A => n3680, B => n8122, C => n3679, D => n8121, Z => 
                           n1201);
   U3784 : AO4 port map( A => n3682, B => n8124, C => n3681, D => n8123, Z => 
                           n1202);
   U3785 : NR4 port map( A => n1204, B => n1205, C => n1206, D => n1207, Z => 
                           n1198);
   U3786 : AO4 port map( A => n3686, B => n8112, C => n3685, D => n8111, Z => 
                           n1204);
   U3787 : AO4 port map( A => n3688, B => n8114, C => n3687, D => n8113, Z => 
                           n1205);
   U3788 : AO4 port map( A => n3690, B => n8116, C => n3689, D => n8115, Z => 
                           n1206);
   U3789 : NR4 port map( A => n1208, B => n1209, C => n1210, D => n1211, Z => 
                           n1197);
   U3790 : AO4 port map( A => n3694, B => n8104, C => n3693, D => n8103, Z => 
                           n1208);
   U3791 : AO4 port map( A => n3696, B => n8106, C => n3695, D => n8105, Z => 
                           n1209);
   U3792 : AO4 port map( A => n3698, B => n8108, C => n3697, D => n8107, Z => 
                           n1210);
   U3793 : NR4 port map( A => n1212, B => n1213, C => n1214, D => n1215, Z => 
                           n1196);
   U3794 : AO4 port map( A => n3702, B => n8096, C => n3701, D => n8095, Z => 
                           n1212);
   U3795 : AO4 port map( A => n3704, B => n8098, C => n3703, D => n8097, Z => 
                           n1213);
   U3796 : AO4 port map( A => n3706, B => n8100, C => n3705, D => n8099, Z => 
                           n1214);
   U3797 : NR4 port map( A => n1220, B => n1221, C => n1222, D => n1223, Z => 
                           n1219);
   U3798 : AO4 port map( A => n3646, B => n8088, C => n3645, D => n8087, Z => 
                           n1220);
   U3799 : AO4 port map( A => n3648, B => n8090, C => n3647, D => n8089, Z => 
                           n1221);
   U3800 : AO4 port map( A => n3650, B => n8092, C => n3649, D => n8091, Z => 
                           n1222);
   U3801 : NR4 port map( A => n1224, B => n1225, C => n1226, D => n1227, Z => 
                           n1218);
   U3802 : AO4 port map( A => n3654, B => n8080, C => n3653, D => n8079, Z => 
                           n1224);
   U3803 : AO4 port map( A => n3656, B => n8082, C => n3655, D => n8081, Z => 
                           n1225);
   U3804 : AO4 port map( A => n3658, B => n8084, C => n3657, D => n8083, Z => 
                           n1226);
   U3805 : NR4 port map( A => n1228, B => n1229, C => n1230, D => n1231, Z => 
                           n1217);
   U3806 : AO4 port map( A => n3662, B => n8072, C => n3661, D => n8071, Z => 
                           n1228);
   U3807 : AO4 port map( A => n3664, B => n8074, C => n3663, D => n8073, Z => 
                           n1229);
   U3808 : AO4 port map( A => n3666, B => n8076, C => n3665, D => n8075, Z => 
                           n1230);
   U3809 : NR4 port map( A => n1232, B => n1233, C => n1234, D => n1235, Z => 
                           n1216);
   U3810 : AO4 port map( A => n3670, B => n8064, C => n3669, D => n8063, Z => 
                           n1232);
   U3811 : AO4 port map( A => n3672, B => n8066, C => n3671, D => n8065, Z => 
                           n1233);
   U3812 : AO4 port map( A => n3674, B => n8068, C => n3673, D => n8067, Z => 
                           n1234);
   U3813 : NR4 port map( A => n1243, B => n1244, C => n1245, D => n1246, Z => 
                           n1242);
   U3814 : AO4 port map( A => n3742, B => n8120, C => n3741, D => n8119, Z => 
                           n1243);
   U3815 : AO4 port map( A => n3744, B => n8122, C => n3743, D => n8121, Z => 
                           n1244);
   U3816 : AO4 port map( A => n3746, B => n8124, C => n3745, D => n8123, Z => 
                           n1245);
   U3817 : NR4 port map( A => n1247, B => n1248, C => n1249, D => n1250, Z => 
                           n1241);
   U3818 : AO4 port map( A => n3750, B => n8112, C => n3749, D => n8111, Z => 
                           n1247);
   U3819 : AO4 port map( A => n3752, B => n8114, C => n3751, D => n8113, Z => 
                           n1248);
   U3820 : AO4 port map( A => n3754, B => n8116, C => n3753, D => n8115, Z => 
                           n1249);
   U3821 : NR4 port map( A => n1251, B => n1252, C => n1253, D => n1254, Z => 
                           n1240);
   U3822 : AO4 port map( A => n3758, B => n8104, C => n3757, D => n8103, Z => 
                           n1251);
   U3823 : AO4 port map( A => n3760, B => n8106, C => n3759, D => n8105, Z => 
                           n1252);
   U3824 : AO4 port map( A => n3762, B => n8108, C => n3761, D => n8107, Z => 
                           n1253);
   U3825 : NR4 port map( A => n1255, B => n1256, C => n1257, D => n1258, Z => 
                           n1239);
   U3826 : AO4 port map( A => n3766, B => n8096, C => n3765, D => n8095, Z => 
                           n1255);
   U3827 : AO4 port map( A => n3768, B => n8098, C => n3767, D => n8097, Z => 
                           n1256);
   U3828 : AO4 port map( A => n3770, B => n8100, C => n3769, D => n8099, Z => 
                           n1257);
   U3829 : NR4 port map( A => n1263, B => n1264, C => n1265, D => n1266, Z => 
                           n1262);
   U3830 : AO4 port map( A => n3710, B => n8088, C => n3709, D => n8087, Z => 
                           n1263);
   U3831 : AO4 port map( A => n3712, B => n8090, C => n3711, D => n8089, Z => 
                           n1264);
   U3832 : AO4 port map( A => n3714, B => n8092, C => n3713, D => n8091, Z => 
                           n1265);
   U3833 : NR4 port map( A => n1267, B => n1268, C => n1269, D => n1270, Z => 
                           n1261);
   U3834 : AO4 port map( A => n3718, B => n8080, C => n3717, D => n8079, Z => 
                           n1267);
   U3835 : AO4 port map( A => n3720, B => n8082, C => n3719, D => n8081, Z => 
                           n1268);
   U3836 : AO4 port map( A => n3722, B => n8084, C => n3721, D => n8083, Z => 
                           n1269);
   U3837 : NR4 port map( A => n1271, B => n1272, C => n1273, D => n1274, Z => 
                           n1260);
   U3838 : AO4 port map( A => n3726, B => n8072, C => n3725, D => n8071, Z => 
                           n1271);
   U3839 : AO4 port map( A => n3728, B => n8074, C => n3727, D => n8073, Z => 
                           n1272);
   U3840 : AO4 port map( A => n3730, B => n8076, C => n3729, D => n8075, Z => 
                           n1273);
   U3841 : NR4 port map( A => n1275, B => n1276, C => n1277, D => n1278, Z => 
                           n1259);
   U3842 : AO4 port map( A => n3734, B => n8064, C => n3733, D => n8063, Z => 
                           n1275);
   U3843 : AO4 port map( A => n3736, B => n8066, C => n3735, D => n8065, Z => 
                           n1276);
   U3844 : AO4 port map( A => n3738, B => n8068, C => n3737, D => n8067, Z => 
                           n1277);
   U3845 : NR4 port map( A => n1287, B => n1288, C => n1289, D => n1290, Z => 
                           n1286);
   U3846 : AO4 port map( A => n3806, B => n8120, C => n3805, D => n8119, Z => 
                           n1287);
   U3847 : AO4 port map( A => n3808, B => n8122, C => n3807, D => n8121, Z => 
                           n1288);
   U3848 : AO4 port map( A => n3810, B => n8124, C => n3809, D => n8123, Z => 
                           n1289);
   U3849 : NR4 port map( A => n1291, B => n1292, C => n1293, D => n1294, Z => 
                           n1285);
   U3850 : AO4 port map( A => n3814, B => n8112, C => n3813, D => n8111, Z => 
                           n1291);
   U3851 : AO4 port map( A => n3816, B => n8114, C => n3815, D => n8113, Z => 
                           n1292);
   U3852 : AO4 port map( A => n3818, B => n8116, C => n3817, D => n8115, Z => 
                           n1293);
   U3853 : NR4 port map( A => n1295, B => n1296, C => n1297, D => n1298, Z => 
                           n1284);
   U3854 : AO4 port map( A => n3822, B => n8104, C => n3821, D => n8103, Z => 
                           n1295);
   U3855 : AO4 port map( A => n3824, B => n8106, C => n3823, D => n8105, Z => 
                           n1296);
   U3856 : AO4 port map( A => n3826, B => n8108, C => n3825, D => n8107, Z => 
                           n1297);
   U3857 : NR4 port map( A => n1299, B => n1300, C => n1301, D => n1302, Z => 
                           n1283);
   U3858 : AO4 port map( A => n3830, B => n8096, C => n3829, D => n8095, Z => 
                           n1299);
   U3859 : AO4 port map( A => n3832, B => n8098, C => n3831, D => n8097, Z => 
                           n1300);
   U3860 : AO4 port map( A => n3834, B => n8100, C => n3833, D => n8099, Z => 
                           n1301);
   U3861 : NR4 port map( A => n1307, B => n1308, C => n1309, D => n1310, Z => 
                           n1306);
   U3862 : AO4 port map( A => n3774, B => n8088, C => n3773, D => n8087, Z => 
                           n1307);
   U3863 : AO4 port map( A => n3776, B => n8090, C => n3775, D => n8089, Z => 
                           n1308);
   U3864 : AO4 port map( A => n3778, B => n8092, C => n3777, D => n8091, Z => 
                           n1309);
   U3865 : NR4 port map( A => n1311, B => n1312, C => n1313, D => n1314, Z => 
                           n1305);
   U3866 : AO4 port map( A => n3782, B => n8080, C => n3781, D => n8079, Z => 
                           n1311);
   U3867 : AO4 port map( A => n3784, B => n8082, C => n3783, D => n8081, Z => 
                           n1312);
   U3868 : AO4 port map( A => n3786, B => n8084, C => n3785, D => n8083, Z => 
                           n1313);
   U3869 : NR4 port map( A => n1315, B => n1316, C => n1317, D => n1318, Z => 
                           n1304);
   U3870 : AO4 port map( A => n3790, B => n8072, C => n3789, D => n8071, Z => 
                           n1315);
   U3871 : AO4 port map( A => n3792, B => n8074, C => n3791, D => n8073, Z => 
                           n1316);
   U3872 : AO4 port map( A => n3794, B => n8076, C => n3793, D => n8075, Z => 
                           n1317);
   U3873 : NR4 port map( A => n1319, B => n1320, C => n1321, D => n1322, Z => 
                           n1303);
   U3874 : AO4 port map( A => n3798, B => n8064, C => n3797, D => n8063, Z => 
                           n1319);
   U3875 : AO4 port map( A => n3800, B => n8066, C => n3799, D => n8065, Z => 
                           n1320);
   U3876 : AO4 port map( A => n3802, B => n8068, C => n3801, D => n8067, Z => 
                           n1321);
   U3877 : NR4 port map( A => n1331, B => n1332, C => n1333, D => n1334, Z => 
                           n1330);
   U3878 : AO4 port map( A => n3870, B => n8120, C => n3869, D => n8119, Z => 
                           n1331);
   U3879 : AO4 port map( A => n3872, B => n8122, C => n3871, D => n8121, Z => 
                           n1332);
   U3880 : AO4 port map( A => n3874, B => n8124, C => n3873, D => n8123, Z => 
                           n1333);
   U3881 : NR4 port map( A => n1335, B => n1336, C => n1337, D => n1338, Z => 
                           n1329);
   U3882 : AO4 port map( A => n3878, B => n8112, C => n3877, D => n8111, Z => 
                           n1335);
   U3883 : AO4 port map( A => n3880, B => n8114, C => n3879, D => n8113, Z => 
                           n1336);
   U3884 : AO4 port map( A => n3882, B => n8116, C => n3881, D => n8115, Z => 
                           n1337);
   U3885 : NR4 port map( A => n1339, B => n1340, C => n1341, D => n1342, Z => 
                           n1328);
   U3886 : AO4 port map( A => n3886, B => n8104, C => n3885, D => n8103, Z => 
                           n1339);
   U3887 : AO4 port map( A => n3888, B => n8106, C => n3887, D => n8105, Z => 
                           n1340);
   U3888 : AO4 port map( A => n3890, B => n8108, C => n3889, D => n8107, Z => 
                           n1341);
   U3889 : NR4 port map( A => n1343, B => n1344, C => n1345, D => n1346, Z => 
                           n1327);
   U3890 : AO4 port map( A => n3894, B => n8096, C => n3893, D => n8095, Z => 
                           n1343);
   U3891 : AO4 port map( A => n3896, B => n8098, C => n3895, D => n8097, Z => 
                           n1344);
   U3892 : AO4 port map( A => n3898, B => n8100, C => n3897, D => n8099, Z => 
                           n1345);
   U3893 : NR4 port map( A => n1351, B => n1352, C => n1353, D => n1354, Z => 
                           n1350);
   U3894 : AO4 port map( A => n3838, B => n8088, C => n3837, D => n8087, Z => 
                           n1351);
   U3895 : AO4 port map( A => n3840, B => n8090, C => n3839, D => n8089, Z => 
                           n1352);
   U3896 : AO4 port map( A => n3842, B => n8092, C => n3841, D => n8091, Z => 
                           n1353);
   U3897 : NR4 port map( A => n1355, B => n1356, C => n1357, D => n1358, Z => 
                           n1349);
   U3898 : AO4 port map( A => n3846, B => n8080, C => n3845, D => n8079, Z => 
                           n1355);
   U3899 : AO4 port map( A => n3848, B => n8082, C => n3847, D => n8081, Z => 
                           n1356);
   U3900 : AO4 port map( A => n3850, B => n8084, C => n3849, D => n8083, Z => 
                           n1357);
   U3901 : NR4 port map( A => n1359, B => n1360, C => n1361, D => n1362, Z => 
                           n1348);
   U3902 : AO4 port map( A => n3854, B => n8072, C => n3853, D => n8071, Z => 
                           n1359);
   U3903 : AO4 port map( A => n3856, B => n8074, C => n3855, D => n8073, Z => 
                           n1360);
   U3904 : AO4 port map( A => n3858, B => n8076, C => n3857, D => n8075, Z => 
                           n1361);
   U3905 : NR4 port map( A => n1363, B => n1364, C => n1365, D => n1366, Z => 
                           n1347);
   U3906 : AO4 port map( A => n3862, B => n8064, C => n3861, D => n8063, Z => 
                           n1363);
   U3907 : AO4 port map( A => n3864, B => n8066, C => n3863, D => n8065, Z => 
                           n1364);
   U3908 : AO4 port map( A => n3866, B => n8068, C => n3865, D => n8067, Z => 
                           n1365);
   U3909 : NR4 port map( A => n1375, B => n1376, C => n1377, D => n1378, Z => 
                           n1374);
   U3910 : AO4 port map( A => n3934, B => n8120, C => n3933, D => n8119, Z => 
                           n1375);
   U3911 : AO4 port map( A => n3936, B => n8122, C => n3935, D => n8121, Z => 
                           n1376);
   U3912 : AO4 port map( A => n3938, B => n8124, C => n3937, D => n8123, Z => 
                           n1377);
   U3913 : NR4 port map( A => n1379, B => n1380, C => n1381, D => n1382, Z => 
                           n1373);
   U3914 : AO4 port map( A => n3942, B => n8112, C => n3941, D => n8111, Z => 
                           n1379);
   U3915 : AO4 port map( A => n3944, B => n8114, C => n3943, D => n8113, Z => 
                           n1380);
   U3916 : AO4 port map( A => n3946, B => n8116, C => n3945, D => n8115, Z => 
                           n1381);
   U3917 : NR4 port map( A => n1383, B => n1384, C => n1385, D => n1386, Z => 
                           n1372);
   U3918 : AO4 port map( A => n3950, B => n8104, C => n3949, D => n8103, Z => 
                           n1383);
   U3919 : AO4 port map( A => n3952, B => n8106, C => n3951, D => n8105, Z => 
                           n1384);
   U3920 : AO4 port map( A => n3954, B => n8108, C => n3953, D => n8107, Z => 
                           n1385);
   U3921 : NR4 port map( A => n1387, B => n1388, C => n1389, D => n1390, Z => 
                           n1371);
   U3922 : AO4 port map( A => n3958, B => n8096, C => n3957, D => n8095, Z => 
                           n1387);
   U3923 : AO4 port map( A => n3960, B => n8098, C => n3959, D => n8097, Z => 
                           n1388);
   U3924 : AO4 port map( A => n3962, B => n8100, C => n3961, D => n8099, Z => 
                           n1389);
   U3925 : NR4 port map( A => n1395, B => n1396, C => n1397, D => n1398, Z => 
                           n1394);
   U3926 : AO4 port map( A => n3902, B => n8088, C => n3901, D => n8087, Z => 
                           n1395);
   U3927 : AO4 port map( A => n3904, B => n8090, C => n3903, D => n8089, Z => 
                           n1396);
   U3928 : AO4 port map( A => n3906, B => n8092, C => n3905, D => n8091, Z => 
                           n1397);
   U3929 : NR4 port map( A => n1399, B => n1400, C => n1401, D => n1402, Z => 
                           n1393);
   U3930 : AO4 port map( A => n3910, B => n8080, C => n3909, D => n8079, Z => 
                           n1399);
   U3931 : AO4 port map( A => n3912, B => n8082, C => n3911, D => n8081, Z => 
                           n1400);
   U3932 : AO4 port map( A => n3914, B => n8084, C => n3913, D => n8083, Z => 
                           n1401);
   U3933 : NR4 port map( A => n1403, B => n1404, C => n1405, D => n1406, Z => 
                           n1392);
   U3934 : AO4 port map( A => n3918, B => n8072, C => n3917, D => n8071, Z => 
                           n1403);
   U3935 : AO4 port map( A => n3920, B => n8074, C => n3919, D => n8073, Z => 
                           n1404);
   U3936 : AO4 port map( A => n3922, B => n8076, C => n3921, D => n8075, Z => 
                           n1405);
   U3937 : NR4 port map( A => n1407, B => n1408, C => n1409, D => n1410, Z => 
                           n1391);
   U3938 : AO4 port map( A => n3926, B => n8064, C => n3925, D => n8063, Z => 
                           n1407);
   U3939 : AO4 port map( A => n3928, B => n8066, C => n3927, D => n8065, Z => 
                           n1408);
   U3940 : AO4 port map( A => n3930, B => n8068, C => n3929, D => n8067, Z => 
                           n1409);
   U3941 : NR4 port map( A => n1418, B => n1419, C => n1420, D => n1421, Z => 
                           n1417);
   U3942 : AO4 port map( A => n3998, B => n8120, C => n3997, D => n8119, Z => 
                           n1418);
   U3943 : AO4 port map( A => n4000, B => n8122, C => n3999, D => n8121, Z => 
                           n1419);
   U3944 : AO4 port map( A => n4002, B => n8124, C => n4001, D => n8123, Z => 
                           n1420);
   U3945 : NR4 port map( A => n1422, B => n1423, C => n1424, D => n1425, Z => 
                           n1416);
   U3946 : AO4 port map( A => n4006, B => n8112, C => n4005, D => n8111, Z => 
                           n1422);
   U3947 : AO4 port map( A => n4008, B => n8114, C => n4007, D => n8113, Z => 
                           n1423);
   U3948 : AO4 port map( A => n4010, B => n8116, C => n4009, D => n8115, Z => 
                           n1424);
   U3949 : NR4 port map( A => n1426, B => n1427, C => n1428, D => n1429, Z => 
                           n1415);
   U3950 : AO4 port map( A => n4014, B => n8104, C => n4013, D => n8103, Z => 
                           n1426);
   U3951 : AO4 port map( A => n4016, B => n8106, C => n4015, D => n8105, Z => 
                           n1427);
   U3952 : AO4 port map( A => n4018, B => n8108, C => n4017, D => n8107, Z => 
                           n1428);
   U3953 : NR4 port map( A => n1430, B => n1431, C => n1432, D => n1433, Z => 
                           n1414);
   U3954 : AO4 port map( A => n4022, B => n8096, C => n4021, D => n8095, Z => 
                           n1430);
   U3955 : AO4 port map( A => n4024, B => n8098, C => n4023, D => n8097, Z => 
                           n1431);
   U3956 : AO4 port map( A => n4026, B => n8100, C => n4025, D => n8099, Z => 
                           n1432);
   U3957 : NR4 port map( A => n1438, B => n1439, C => n1440, D => n1441, Z => 
                           n1437);
   U3958 : AO4 port map( A => n3966, B => n8088, C => n3965, D => n8087, Z => 
                           n1438);
   U3959 : AO4 port map( A => n3968, B => n8090, C => n3967, D => n8089, Z => 
                           n1439);
   U3960 : AO4 port map( A => n3970, B => n8092, C => n3969, D => n8091, Z => 
                           n1440);
   U3961 : NR4 port map( A => n1442, B => n1443, C => n1444, D => n1445, Z => 
                           n1436);
   U3962 : AO4 port map( A => n3974, B => n8080, C => n3973, D => n8079, Z => 
                           n1442);
   U3963 : AO4 port map( A => n3976, B => n8082, C => n3975, D => n8081, Z => 
                           n1443);
   U3964 : AO4 port map( A => n3978, B => n8084, C => n3977, D => n8083, Z => 
                           n1444);
   U3965 : NR4 port map( A => n1446, B => n1447, C => n1448, D => n1449, Z => 
                           n1435);
   U3966 : AO4 port map( A => n3982, B => n8072, C => n3981, D => n8071, Z => 
                           n1446);
   U3967 : AO4 port map( A => n3984, B => n8074, C => n3983, D => n8073, Z => 
                           n1447);
   U3968 : AO4 port map( A => n3986, B => n8076, C => n3985, D => n8075, Z => 
                           n1448);
   U3969 : NR4 port map( A => n1450, B => n1451, C => n1452, D => n1453, Z => 
                           n1434);
   U3970 : AO4 port map( A => n3990, B => n8064, C => n3989, D => n8063, Z => 
                           n1450);
   U3971 : AO4 port map( A => n3992, B => n8066, C => n3991, D => n8065, Z => 
                           n1451);
   U3972 : AO4 port map( A => n3994, B => n8068, C => n3993, D => n8067, Z => 
                           n1452);
   U3973 : NR4 port map( A => n1462, B => n1463, C => n1464, D => n1465, Z => 
                           n1461);
   U3974 : AO4 port map( A => n4062, B => n8120, C => n4061, D => n8119, Z => 
                           n1462);
   U3975 : AO4 port map( A => n4064, B => n8122, C => n4063, D => n8121, Z => 
                           n1463);
   U3976 : AO4 port map( A => n4066, B => n8124, C => n4065, D => n8123, Z => 
                           n1464);
   U3977 : NR4 port map( A => n1466, B => n1467, C => n1468, D => n1469, Z => 
                           n1460);
   U3978 : AO4 port map( A => n4070, B => n8112, C => n4069, D => n8111, Z => 
                           n1466);
   U3979 : AO4 port map( A => n4072, B => n8114, C => n4071, D => n8113, Z => 
                           n1467);
   U3980 : AO4 port map( A => n4074, B => n8116, C => n4073, D => n8115, Z => 
                           n1468);
   U3981 : NR4 port map( A => n1470, B => n1471, C => n1472, D => n1473, Z => 
                           n1459);
   U3982 : AO4 port map( A => n4078, B => n8104, C => n4077, D => n8103, Z => 
                           n1470);
   U3983 : AO4 port map( A => n4080, B => n8106, C => n4079, D => n8105, Z => 
                           n1471);
   U3984 : AO4 port map( A => n4082, B => n8108, C => n4081, D => n8107, Z => 
                           n1472);
   U3985 : NR4 port map( A => n1474, B => n1475, C => n1476, D => n1477, Z => 
                           n1458);
   U3986 : AO4 port map( A => n4086, B => n8096, C => n4085, D => n8095, Z => 
                           n1474);
   U3987 : AO4 port map( A => n4088, B => n8098, C => n4087, D => n8097, Z => 
                           n1475);
   U3988 : AO4 port map( A => n4090, B => n8100, C => n4089, D => n8099, Z => 
                           n1476);
   U3989 : NR4 port map( A => n1482, B => n1483, C => n1484, D => n1485, Z => 
                           n1481);
   U3990 : AO4 port map( A => n4030, B => n8088, C => n4029, D => n8087, Z => 
                           n1482);
   U3991 : AO4 port map( A => n4032, B => n8090, C => n4031, D => n8089, Z => 
                           n1483);
   U3992 : AO4 port map( A => n4034, B => n8092, C => n4033, D => n8091, Z => 
                           n1484);
   U3993 : NR4 port map( A => n1486, B => n1487, C => n1488, D => n1489, Z => 
                           n1480);
   U3994 : AO4 port map( A => n4038, B => n8080, C => n4037, D => n8079, Z => 
                           n1486);
   U3995 : AO4 port map( A => n4040, B => n8082, C => n4039, D => n8081, Z => 
                           n1487);
   U3996 : AO4 port map( A => n4042, B => n8084, C => n4041, D => n8083, Z => 
                           n1488);
   U3997 : NR4 port map( A => n1490, B => n1491, C => n1492, D => n1493, Z => 
                           n1479);
   U3998 : AO4 port map( A => n4046, B => n8072, C => n4045, D => n8071, Z => 
                           n1490);
   U3999 : AO4 port map( A => n4048, B => n8074, C => n4047, D => n8073, Z => 
                           n1491);
   U4000 : AO4 port map( A => n4050, B => n8076, C => n4049, D => n8075, Z => 
                           n1492);
   U4001 : NR4 port map( A => n1494, B => n1495, C => n1496, D => n1497, Z => 
                           n1478);
   U4002 : AO4 port map( A => n4054, B => n8064, C => n4053, D => n8063, Z => 
                           n1494);
   U4003 : AO4 port map( A => n4056, B => n8066, C => n4055, D => n8065, Z => 
                           n1495);
   U4004 : AO4 port map( A => n4058, B => n8068, C => n4057, D => n8067, Z => 
                           n1496);
   U4005 : NR4 port map( A => n1506, B => n1507, C => n1508, D => n1509, Z => 
                           n1505);
   U4006 : AO4 port map( A => n4126, B => n8120, C => n4125, D => n8119, Z => 
                           n1506);
   U4007 : AO4 port map( A => n4128, B => n8122, C => n4127, D => n8121, Z => 
                           n1507);
   U4008 : AO4 port map( A => n4130, B => n8124, C => n4129, D => n8123, Z => 
                           n1508);
   U4009 : NR4 port map( A => n1510, B => n1511, C => n1512, D => n1513, Z => 
                           n1504);
   U4010 : AO4 port map( A => n4134, B => n8112, C => n4133, D => n8111, Z => 
                           n1510);
   U4011 : AO4 port map( A => n4136, B => n8114, C => n4135, D => n8113, Z => 
                           n1511);
   U4012 : AO4 port map( A => n4138, B => n8116, C => n4137, D => n8115, Z => 
                           n1512);
   U4013 : NR4 port map( A => n1514, B => n1515, C => n1516, D => n1517, Z => 
                           n1503);
   U4014 : AO4 port map( A => n4142, B => n8104, C => n4141, D => n8103, Z => 
                           n1514);
   U4015 : AO4 port map( A => n4144, B => n8106, C => n4143, D => n8105, Z => 
                           n1515);
   U4016 : AO4 port map( A => n4146, B => n8108, C => n4145, D => n8107, Z => 
                           n1516);
   U4017 : NR4 port map( A => n1518, B => n1519, C => n1520, D => n1521, Z => 
                           n1502);
   U4018 : AO4 port map( A => n4150, B => n8096, C => n4149, D => n8095, Z => 
                           n1518);
   U4019 : AO4 port map( A => n4152, B => n8098, C => n4151, D => n8097, Z => 
                           n1519);
   U4020 : AO4 port map( A => n4154, B => n8100, C => n4153, D => n8099, Z => 
                           n1520);
   U4021 : NR4 port map( A => n1526, B => n1527, C => n1528, D => n1529, Z => 
                           n1525);
   U4022 : AO4 port map( A => n4094, B => n8088, C => n4093, D => n8087, Z => 
                           n1526);
   U4023 : AO4 port map( A => n4096, B => n8090, C => n4095, D => n8089, Z => 
                           n1527);
   U4024 : AO4 port map( A => n4098, B => n8092, C => n4097, D => n8091, Z => 
                           n1528);
   U4025 : NR4 port map( A => n1530, B => n1531, C => n1532, D => n1533, Z => 
                           n1524);
   U4026 : AO4 port map( A => n4102, B => n8080, C => n4101, D => n8079, Z => 
                           n1530);
   U4027 : AO4 port map( A => n4104, B => n8082, C => n4103, D => n8081, Z => 
                           n1531);
   U4028 : AO4 port map( A => n4106, B => n8084, C => n4105, D => n8083, Z => 
                           n1532);
   U4029 : NR4 port map( A => n1534, B => n1535, C => n1536, D => n1537, Z => 
                           n1523);
   U4030 : AO4 port map( A => n4110, B => n8072, C => n4109, D => n8071, Z => 
                           n1534);
   U4031 : AO4 port map( A => n4112, B => n8074, C => n4111, D => n8073, Z => 
                           n1535);
   U4032 : AO4 port map( A => n4114, B => n8076, C => n4113, D => n8075, Z => 
                           n1536);
   U4033 : NR4 port map( A => n1538, B => n1539, C => n1540, D => n1541, Z => 
                           n1522);
   U4034 : AO4 port map( A => n4118, B => n8064, C => n4117, D => n8063, Z => 
                           n1538);
   U4035 : AO4 port map( A => n4120, B => n8066, C => n4119, D => n8065, Z => 
                           n1539);
   U4036 : AO4 port map( A => n4122, B => n8068, C => n4121, D => n8067, Z => 
                           n1540);
   U4037 : NR4 port map( A => n1550, B => n1551, C => n1552, D => n1553, Z => 
                           n1549);
   U4038 : AO4 port map( A => n4190, B => n8120, C => n4189, D => n8119, Z => 
                           n1550);
   U4039 : AO4 port map( A => n4192, B => n8122, C => n4191, D => n8121, Z => 
                           n1551);
   U4040 : AO4 port map( A => n4194, B => n8124, C => n4193, D => n8123, Z => 
                           n1552);
   U4041 : NR4 port map( A => n1554, B => n1555, C => n1556, D => n1557, Z => 
                           n1548);
   U4042 : AO4 port map( A => n4198, B => n8112, C => n4197, D => n8111, Z => 
                           n1554);
   U4043 : AO4 port map( A => n4200, B => n8114, C => n4199, D => n8113, Z => 
                           n1555);
   U4044 : AO4 port map( A => n4202, B => n8116, C => n4201, D => n8115, Z => 
                           n1556);
   U4045 : NR4 port map( A => n1558, B => n1559, C => n1560, D => n1561, Z => 
                           n1547);
   U4046 : AO4 port map( A => n4206, B => n8104, C => n4205, D => n8103, Z => 
                           n1558);
   U4047 : AO4 port map( A => n4208, B => n8106, C => n4207, D => n8105, Z => 
                           n1559);
   U4048 : AO4 port map( A => n4210, B => n8108, C => n4209, D => n8107, Z => 
                           n1560);
   U4049 : NR4 port map( A => n1562, B => n1563, C => n1564, D => n1565, Z => 
                           n1546);
   U4050 : AO4 port map( A => n4214, B => n8096, C => n4213, D => n8095, Z => 
                           n1562);
   U4051 : AO4 port map( A => n4216, B => n8098, C => n4215, D => n8097, Z => 
                           n1563);
   U4052 : AO4 port map( A => n4218, B => n8100, C => n4217, D => n8099, Z => 
                           n1564);
   U4053 : NR4 port map( A => n1570, B => n1571, C => n1572, D => n1573, Z => 
                           n1569);
   U4054 : AO4 port map( A => n4158, B => n8088, C => n4157, D => n8087, Z => 
                           n1570);
   U4055 : AO4 port map( A => n4160, B => n8090, C => n4159, D => n8089, Z => 
                           n1571);
   U4056 : AO4 port map( A => n4162, B => n8092, C => n4161, D => n8091, Z => 
                           n1572);
   U4057 : NR4 port map( A => n1574, B => n1575, C => n1576, D => n1577, Z => 
                           n1568);
   U4058 : AO4 port map( A => n4166, B => n8080, C => n4165, D => n8079, Z => 
                           n1574);
   U4059 : AO4 port map( A => n4168, B => n8082, C => n4167, D => n8081, Z => 
                           n1575);
   U4060 : AO4 port map( A => n4170, B => n8084, C => n4169, D => n8083, Z => 
                           n1576);
   U4061 : NR4 port map( A => n1578, B => n1579, C => n1580, D => n1581, Z => 
                           n1567);
   U4062 : AO4 port map( A => n4174, B => n8072, C => n4173, D => n8071, Z => 
                           n1578);
   U4063 : AO4 port map( A => n4176, B => n8074, C => n4175, D => n8073, Z => 
                           n1579);
   U4064 : AO4 port map( A => n4178, B => n8076, C => n4177, D => n8075, Z => 
                           n1580);
   U4065 : NR4 port map( A => n1582, B => n1583, C => n1584, D => n1585, Z => 
                           n1566);
   U4066 : AO4 port map( A => n4182, B => n8064, C => n4181, D => n8063, Z => 
                           n1582);
   U4067 : AO4 port map( A => n4184, B => n8066, C => n4183, D => n8065, Z => 
                           n1583);
   U4068 : AO4 port map( A => n4186, B => n8068, C => n4185, D => n8067, Z => 
                           n1584);
   U4069 : NR4 port map( A => n1594, B => n1595, C => n1596, D => n1597, Z => 
                           n1593);
   U4070 : AO4 port map( A => n4254, B => n8120, C => n4253, D => n8119, Z => 
                           n1594);
   U4071 : AO4 port map( A => n4256, B => n8122, C => n4255, D => n8121, Z => 
                           n1595);
   U4072 : AO4 port map( A => n4258, B => n8124, C => n4257, D => n8123, Z => 
                           n1596);
   U4073 : NR4 port map( A => n1598, B => n1599, C => n1600, D => n1601, Z => 
                           n1592);
   U4074 : AO4 port map( A => n4262, B => n8112, C => n4261, D => n8111, Z => 
                           n1598);
   U4075 : AO4 port map( A => n4264, B => n8114, C => n4263, D => n8113, Z => 
                           n1599);
   U4076 : AO4 port map( A => n4266, B => n8116, C => n4265, D => n8115, Z => 
                           n1600);
   U4077 : NR4 port map( A => n1602, B => n1603, C => n1604, D => n1605, Z => 
                           n1591);
   U4078 : AO4 port map( A => n4270, B => n8104, C => n4269, D => n8103, Z => 
                           n1602);
   U4079 : AO4 port map( A => n4272, B => n8106, C => n4271, D => n8105, Z => 
                           n1603);
   U4080 : AO4 port map( A => n4274, B => n8108, C => n4273, D => n8107, Z => 
                           n1604);
   U4081 : NR4 port map( A => n1606, B => n1607, C => n1608, D => n1609, Z => 
                           n1590);
   U4082 : AO4 port map( A => n4278, B => n8096, C => n4277, D => n8095, Z => 
                           n1606);
   U4083 : AO4 port map( A => n4280, B => n8098, C => n4279, D => n8097, Z => 
                           n1607);
   U4084 : AO4 port map( A => n4282, B => n8100, C => n4281, D => n8099, Z => 
                           n1608);
   U4085 : NR4 port map( A => n1614, B => n1615, C => n1616, D => n1617, Z => 
                           n1613);
   U4086 : AO4 port map( A => n4222, B => n8088, C => n4221, D => n8087, Z => 
                           n1614);
   U4087 : AO4 port map( A => n4224, B => n8090, C => n4223, D => n8089, Z => 
                           n1615);
   U4088 : AO4 port map( A => n4226, B => n8092, C => n4225, D => n8091, Z => 
                           n1616);
   U4089 : NR4 port map( A => n1618, B => n1619, C => n1620, D => n1621, Z => 
                           n1612);
   U4090 : AO4 port map( A => n4230, B => n8080, C => n4229, D => n8079, Z => 
                           n1618);
   U4091 : AO4 port map( A => n4232, B => n8082, C => n4231, D => n8081, Z => 
                           n1619);
   U4092 : AO4 port map( A => n4234, B => n8084, C => n4233, D => n8083, Z => 
                           n1620);
   U4093 : NR4 port map( A => n1622, B => n1623, C => n1624, D => n1625, Z => 
                           n1611);
   U4094 : AO4 port map( A => n4238, B => n8072, C => n4237, D => n8071, Z => 
                           n1622);
   U4095 : AO4 port map( A => n4240, B => n8074, C => n4239, D => n8073, Z => 
                           n1623);
   U4096 : AO4 port map( A => n4242, B => n8076, C => n4241, D => n8075, Z => 
                           n1624);
   U4097 : NR4 port map( A => n1626, B => n1627, C => n1628, D => n1629, Z => 
                           n1610);
   U4098 : AO4 port map( A => n4246, B => n8064, C => n4245, D => n8063, Z => 
                           n1626);
   U4099 : AO4 port map( A => n4248, B => n8066, C => n4247, D => n8065, Z => 
                           n1627);
   U4100 : AO4 port map( A => n4250, B => n8068, C => n4249, D => n8067, Z => 
                           n1628);
   U4101 : NR4 port map( A => n1638, B => n1639, C => n1640, D => n1641, Z => 
                           n1637);
   U4102 : AO4 port map( A => n4319, B => n8120, C => n4318, D => n8119, Z => 
                           n1638);
   U4103 : AO4 port map( A => n4321, B => n8122, C => n4320, D => n8121, Z => 
                           n1639);
   U4104 : AO4 port map( A => n4323, B => n8124, C => n4322, D => n8123, Z => 
                           n1640);
   U4105 : NR4 port map( A => n1642, B => n1643, C => n1644, D => n1645, Z => 
                           n1636);
   U4106 : AO4 port map( A => n4327, B => n8112, C => n4326, D => n8111, Z => 
                           n1642);
   U4107 : AO4 port map( A => n4329, B => n8114, C => n4328, D => n8113, Z => 
                           n1643);
   U4108 : AO4 port map( A => n4331, B => n8116, C => n4330, D => n8115, Z => 
                           n1644);
   U4109 : NR4 port map( A => n1646, B => n1647, C => n1648, D => n1649, Z => 
                           n1635);
   U4110 : AO4 port map( A => n4335, B => n8104, C => n4334, D => n8103, Z => 
                           n1646);
   U4111 : AO4 port map( A => n4337, B => n8106, C => n4336, D => n8105, Z => 
                           n1647);
   U4112 : AO4 port map( A => n4339, B => n8108, C => n4338, D => n8107, Z => 
                           n1648);
   U4113 : NR4 port map( A => n1650, B => n1651, C => n1652, D => n1653, Z => 
                           n1634);
   U4114 : AO4 port map( A => n4343, B => n8096, C => n4342, D => n8095, Z => 
                           n1650);
   U4115 : AO4 port map( A => n4345, B => n8098, C => n4344, D => n8097, Z => 
                           n1651);
   U4116 : AO4 port map( A => n4347, B => n8100, C => n4346, D => n8099, Z => 
                           n1652);
   U4117 : NR4 port map( A => n1658, B => n1659, C => n1660, D => n1661, Z => 
                           n1657);
   U4118 : AO4 port map( A => n4287, B => n8088, C => n4286, D => n8087, Z => 
                           n1658);
   U4119 : AO4 port map( A => n4289, B => n8090, C => n4288, D => n8089, Z => 
                           n1659);
   U4120 : AO4 port map( A => n4291, B => n8092, C => n4290, D => n8091, Z => 
                           n1660);
   U4121 : NR4 port map( A => n1662, B => n1663, C => n1664, D => n1665, Z => 
                           n1656);
   U4122 : AO4 port map( A => n4295, B => n8080, C => n4294, D => n8079, Z => 
                           n1662);
   U4123 : AO4 port map( A => n4297, B => n8082, C => n4296, D => n8081, Z => 
                           n1663);
   U4124 : AO4 port map( A => n4299, B => n8084, C => n4298, D => n8083, Z => 
                           n1664);
   U4125 : NR4 port map( A => n1666, B => n1667, C => n1668, D => n1669, Z => 
                           n1655);
   U4126 : AO4 port map( A => n4303, B => n8072, C => n4302, D => n8071, Z => 
                           n1666);
   U4127 : AO4 port map( A => n4305, B => n8074, C => n4304, D => n8073, Z => 
                           n1667);
   U4128 : AO4 port map( A => n4307, B => n8076, C => n4306, D => n8075, Z => 
                           n1668);
   U4129 : NR4 port map( A => n1670, B => n1671, C => n1672, D => n1673, Z => 
                           n1654);
   U4130 : AO4 port map( A => n4311, B => n8064, C => n4310, D => n8063, Z => 
                           n1670);
   U4131 : AO4 port map( A => n4313, B => n8066, C => n4312, D => n8065, Z => 
                           n1671);
   U4132 : AO4 port map( A => n4315, B => n8068, C => n4314, D => n8067, Z => 
                           n1672);
   U4133 : NR4 port map( A => n1682, B => n1683, C => n1684, D => n1685, Z => 
                           n1681);
   U4134 : AO4 port map( A => n4383, B => n8120, C => n4382, D => n8119, Z => 
                           n1682);
   U4135 : AO4 port map( A => n4385, B => n8122, C => n4384, D => n8121, Z => 
                           n1683);
   U4136 : AO4 port map( A => n4387, B => n8124, C => n4386, D => n8123, Z => 
                           n1684);
   U4137 : NR4 port map( A => n1686, B => n1687, C => n1688, D => n1689, Z => 
                           n1680);
   U4138 : AO4 port map( A => n4391, B => n8112, C => n4390, D => n8111, Z => 
                           n1686);
   U4139 : AO4 port map( A => n4393, B => n8114, C => n4392, D => n8113, Z => 
                           n1687);
   U4140 : AO4 port map( A => n4395, B => n8116, C => n4394, D => n8115, Z => 
                           n1688);
   U4141 : NR4 port map( A => n1690, B => n1691, C => n1692, D => n1693, Z => 
                           n1679);
   U4142 : AO4 port map( A => n4399, B => n8104, C => n4398, D => n8103, Z => 
                           n1690);
   U4143 : AO4 port map( A => n4401, B => n8106, C => n4400, D => n8105, Z => 
                           n1691);
   U4144 : AO4 port map( A => n4403, B => n8108, C => n4402, D => n8107, Z => 
                           n1692);
   U4145 : NR4 port map( A => n1694, B => n1695, C => n1696, D => n1697, Z => 
                           n1678);
   U4146 : AO4 port map( A => n4407, B => n8096, C => n4406, D => n8095, Z => 
                           n1694);
   U4147 : AO4 port map( A => n4409, B => n8098, C => n4408, D => n8097, Z => 
                           n1695);
   U4148 : AO4 port map( A => n4411, B => n8100, C => n4410, D => n8099, Z => 
                           n1696);
   U4149 : NR4 port map( A => n1702, B => n1703, C => n1704, D => n1705, Z => 
                           n1701);
   U4150 : AO4 port map( A => n4351, B => n8088, C => n4350, D => n8087, Z => 
                           n1702);
   U4151 : AO4 port map( A => n4353, B => n8090, C => n4352, D => n8089, Z => 
                           n1703);
   U4152 : AO4 port map( A => n4355, B => n8092, C => n4354, D => n8091, Z => 
                           n1704);
   U4153 : NR4 port map( A => n1706, B => n1707, C => n1708, D => n1709, Z => 
                           n1700);
   U4154 : AO4 port map( A => n4359, B => n8080, C => n4358, D => n8079, Z => 
                           n1706);
   U4155 : AO4 port map( A => n4361, B => n8082, C => n4360, D => n8081, Z => 
                           n1707);
   U4156 : AO4 port map( A => n4363, B => n8084, C => n4362, D => n8083, Z => 
                           n1708);
   U4157 : NR4 port map( A => n1710, B => n1711, C => n1712, D => n1713, Z => 
                           n1699);
   U4158 : AO4 port map( A => n4367, B => n8072, C => n4366, D => n8071, Z => 
                           n1710);
   U4159 : AO4 port map( A => n4369, B => n8074, C => n4368, D => n8073, Z => 
                           n1711);
   U4160 : AO4 port map( A => n4371, B => n8076, C => n4370, D => n8075, Z => 
                           n1712);
   U4161 : NR4 port map( A => n1714, B => n1715, C => n1716, D => n1717, Z => 
                           n1698);
   U4162 : AO4 port map( A => n4375, B => n8064, C => n4374, D => n8063, Z => 
                           n1714);
   U4163 : AO4 port map( A => n4377, B => n8066, C => n4376, D => n8065, Z => 
                           n1715);
   U4164 : AO4 port map( A => n4379, B => n8068, C => n4378, D => n8067, Z => 
                           n1716);
   U4165 : NR4 port map( A => n1726, B => n1727, C => n1728, D => n1729, Z => 
                           n1725);
   U4166 : AO4 port map( A => n4447, B => n8120, C => n4446, D => n8119, Z => 
                           n1726);
   U4167 : AO4 port map( A => n4449, B => n8122, C => n4448, D => n8121, Z => 
                           n1727);
   U4168 : AO4 port map( A => n4451, B => n8124, C => n4450, D => n8123, Z => 
                           n1728);
   U4169 : NR4 port map( A => n1730, B => n1731, C => n1732, D => n1733, Z => 
                           n1724);
   U4170 : AO4 port map( A => n4455, B => n8112, C => n4454, D => n8111, Z => 
                           n1730);
   U4171 : AO4 port map( A => n4457, B => n8114, C => n4456, D => n8113, Z => 
                           n1731);
   U4172 : AO4 port map( A => n4459, B => n8116, C => n4458, D => n8115, Z => 
                           n1732);
   U4173 : NR4 port map( A => n1734, B => n1735, C => n1736, D => n1737, Z => 
                           n1723);
   U4174 : AO4 port map( A => n4463, B => n8104, C => n4462, D => n8103, Z => 
                           n1734);
   U4175 : AO4 port map( A => n4465, B => n8106, C => n4464, D => n8105, Z => 
                           n1735);
   U4176 : AO4 port map( A => n4467, B => n8108, C => n4466, D => n8107, Z => 
                           n1736);
   U4177 : NR4 port map( A => n1738, B => n1739, C => n1740, D => n1741, Z => 
                           n1722);
   U4178 : AO4 port map( A => n4471, B => n8096, C => n4470, D => n8095, Z => 
                           n1738);
   U4179 : AO4 port map( A => n4473, B => n8098, C => n4472, D => n8097, Z => 
                           n1739);
   U4180 : AO4 port map( A => n4475, B => n8100, C => n4474, D => n8099, Z => 
                           n1740);
   U4181 : NR4 port map( A => n1746, B => n1747, C => n1748_port, D => 
                           n1749_port, Z => n1745);
   U4182 : AO4 port map( A => n4415, B => n8088, C => n4414, D => n8087, Z => 
                           n1746);
   U4183 : AO4 port map( A => n4417, B => n8090, C => n4416, D => n8089, Z => 
                           n1747);
   U4184 : AO4 port map( A => n4419, B => n8092, C => n4418, D => n8091, Z => 
                           n1748_port);
   U4185 : NR4 port map( A => n1750_port, B => n1751_port, C => n1752_port, D 
                           => n1753_port, Z => n1744);
   U4186 : AO4 port map( A => n4423, B => n8080, C => n4422, D => n8079, Z => 
                           n1750_port);
   U4187 : AO4 port map( A => n4425, B => n8082, C => n4424, D => n8081, Z => 
                           n1751_port);
   U4188 : AO4 port map( A => n4427, B => n8084, C => n4426, D => n8083, Z => 
                           n1752_port);
   U4189 : NR4 port map( A => n1754_port, B => n1755, C => n1756, D => n1757, Z
                           => n1743);
   U4190 : AO4 port map( A => n4431, B => n8072, C => n4430, D => n8071, Z => 
                           n1754_port);
   U4191 : AO4 port map( A => n4433, B => n8074, C => n4432, D => n8073, Z => 
                           n1755);
   U4192 : AO4 port map( A => n4435, B => n8076, C => n4434, D => n8075, Z => 
                           n1756);
   U4193 : NR4 port map( A => n1758, B => n1759, C => n1760, D => n1761, Z => 
                           n1742);
   U4194 : AO4 port map( A => n4439, B => n8064, C => n4438, D => n8063, Z => 
                           n1758);
   U4195 : AO4 port map( A => n4441, B => n8066, C => n4440, D => n8065, Z => 
                           n1759);
   U4196 : AO4 port map( A => n4443, B => n8068, C => n4442, D => n8067, Z => 
                           n1760);
   U4197 : NR4 port map( A => n1769, B => n1770, C => n1771, D => n1772, Z => 
                           n1768);
   U4198 : AO4 port map( A => n4511, B => n8120, C => n4510, D => n8119, Z => 
                           n1769);
   U4199 : AO4 port map( A => n4513, B => n8122, C => n4512, D => n8121, Z => 
                           n1770);
   U4200 : AO4 port map( A => n4515, B => n8124, C => n4514, D => n8123, Z => 
                           n1771);
   U4201 : NR4 port map( A => n1782, B => n1783, C => n1784, D => n1785, Z => 
                           n1767);
   U4202 : AO4 port map( A => n4519, B => n8112, C => n4518, D => n8111, Z => 
                           n1782);
   U4203 : AO4 port map( A => n4521, B => n8114, C => n4520, D => n8113, Z => 
                           n1783);
   U4204 : AO4 port map( A => n4523, B => n8116, C => n4522, D => n8115, Z => 
                           n1784);
   U4205 : NR4 port map( A => n1792, B => n1793, C => n1794, D => n1795, Z => 
                           n1766);
   U4206 : AO4 port map( A => n4527, B => n8104, C => n4526, D => n8103, Z => 
                           n1792);
   U4207 : AO4 port map( A => n4529, B => n8106, C => n4528, D => n8105, Z => 
                           n1793);
   U4208 : AO4 port map( A => n4531, B => n8108, C => n4530, D => n8107, Z => 
                           n1794);
   U4209 : NR4 port map( A => n1799, B => n1800, C => n1801, D => n1802, Z => 
                           n1765);
   U4210 : AO4 port map( A => n4535, B => n8096, C => n4534, D => n8095, Z => 
                           n1799);
   U4211 : AO4 port map( A => n4537, B => n8098, C => n4536, D => n8097, Z => 
                           n1800);
   U4212 : AO4 port map( A => n4539, B => n8100, C => n4538, D => n8099, Z => 
                           n1801);
   U4213 : NR4 port map( A => n1811, B => n1812, C => n1813, D => n1814, Z => 
                           n1810);
   U4214 : AO4 port map( A => n4479, B => n8088, C => n4478, D => n8087, Z => 
                           n1811);
   U4215 : AO4 port map( A => n4481, B => n8090, C => n4480, D => n8089, Z => 
                           n1812);
   U4216 : AO4 port map( A => n4483, B => n8092, C => n4482, D => n8091, Z => 
                           n1813);
   U4217 : NR4 port map( A => n1818, B => n1819, C => n1820, D => n1821, Z => 
                           n1809);
   U4218 : AO4 port map( A => n4487, B => n8080, C => n4486, D => n8079, Z => 
                           n1818);
   U4219 : AO4 port map( A => n4489, B => n8082, C => n4488, D => n8081, Z => 
                           n1819);
   U4220 : AO4 port map( A => n4491, B => n8084, C => n4490, D => n8083, Z => 
                           n1820);
   U4221 : NR4 port map( A => n1824, B => n1825, C => n1826, D => n1827, Z => 
                           n1808);
   U4222 : AO4 port map( A => n4495, B => n8072, C => n4494, D => n8071, Z => 
                           n1824);
   U4223 : AO4 port map( A => n4497, B => n8074, C => n4496, D => n8073, Z => 
                           n1825);
   U4224 : AO4 port map( A => n4499, B => n8076, C => n4498, D => n8075, Z => 
                           n1826);
   U4225 : NR4 port map( A => n1835, B => n1836, C => n1837, D => n1838, Z => 
                           n1807);
   U4226 : AO4 port map( A => n4503, B => n8064, C => n4502, D => n8063, Z => 
                           n1835);
   U4227 : AO4 port map( A => n4505, B => n8066, C => n4504, D => n8065, Z => 
                           n1836);
   U4228 : AO4 port map( A => n4507, B => n8068, C => n4506, D => n8067, Z => 
                           n1837);
   U4229 : EON1 port map( A => KEY_NUMB_I(1), B => n8302, C => n8302, D => 
                           n6648, Z => n1844);
   U4230 : EON1 port map( A => KEY_NUMB_I(0), B => n8302, C => n8302, D => 
                           n6649, Z => n1843);
   U4231 : EON1 port map( A => KEY_NUMB_I(2), B => n8302, C => n8302, D => 
                           n6647, Z => n1833);
   U4232 : EON1 port map( A => KEY_NUMB_I(3), B => n8302, C => n8302, D => 
                           n6646, Z => n1834);
   U4233 : EON1 port map( A => KEY_NUMB_I(5), B => n8302, C => n8302, D => 
                           n6644, Z => n1806);
   U4234 : EON1 port map( A => KEY_NUMB_I(4), B => n8302, C => n8302, D => 
                           n6645, Z => n1805);
   U4235 : IVI port map( A => GET_KEY_I, Z => n8302);
   U4236 : AO4 port map( A => n2531, B => n8126, C => n2530, D => n8125, Z => 
                           n350);
   U4237 : AO4 port map( A => n2539, B => n8118, C => n2538, D => n8117, Z => 
                           n362);
   U4238 : AO4 port map( A => n2547, B => n8110, C => n2546, D => n8109, Z => 
                           n374);
   U4239 : AO4 port map( A => n2555, B => n8102, C => n2554, D => n8101, Z => 
                           n386);
   U4240 : AO4 port map( A => n2499, B => n8094, C => n2498, D => n8093, Z => 
                           n402);
   U4241 : AO4 port map( A => n2507, B => n8086, C => n2506, D => n8085, Z => 
                           n414);
   U4242 : AO4 port map( A => n2515, B => n8078, C => n2514, D => n8077, Z => 
                           n426);
   U4243 : AO4 port map( A => n2523, B => n8070, C => n2522, D => n8069, Z => 
                           n438);
   U4244 : AO4 port map( A => n2595, B => n8126, C => n2594, D => n8125, Z => 
                           n458);
   U4245 : AO4 port map( A => n2603, B => n8118, C => n2602, D => n8117, Z => 
                           n462);
   U4246 : AO4 port map( A => n2611, B => n8110, C => n2610, D => n8109, Z => 
                           n466);
   U4247 : AO4 port map( A => n2619, B => n8102, C => n2618, D => n8101, Z => 
                           n470);
   U4248 : AO4 port map( A => n2563, B => n8094, C => n2562, D => n8093, Z => 
                           n478);
   U4249 : AO4 port map( A => n2571, B => n8086, C => n2570, D => n8085, Z => 
                           n482);
   U4250 : AO4 port map( A => n2579, B => n8078, C => n2578, D => n8077, Z => 
                           n486);
   U4251 : AO4 port map( A => n2587, B => n8070, C => n2586, D => n8069, Z => 
                           n490);
   U4252 : AO4 port map( A => n2659, B => n8126, C => n2658, D => n8125, Z => 
                           n502);
   U4253 : AO4 port map( A => n2667, B => n8118, C => n2666, D => n8117, Z => 
                           n506);
   U4254 : AO4 port map( A => n2675, B => n8110, C => n2674, D => n8109, Z => 
                           n510);
   U4255 : AO4 port map( A => n2683, B => n8102, C => n2682, D => n8101, Z => 
                           n514);
   U4256 : AO4 port map( A => n2627, B => n8094, C => n2626, D => n8093, Z => 
                           n522);
   U4257 : AO4 port map( A => n2635, B => n8086, C => n2634, D => n8085, Z => 
                           n526);
   U4258 : AO4 port map( A => n2643, B => n8078, C => n2642, D => n8077, Z => 
                           n530);
   U4259 : AO4 port map( A => n2651, B => n8070, C => n2650, D => n8069, Z => 
                           n534);
   U4260 : AO4 port map( A => n2723, B => n8126, C => n2722, D => n8125, Z => 
                           n546);
   U4261 : AO4 port map( A => n2731, B => n8118, C => n2730, D => n8117, Z => 
                           n550);
   U4262 : AO4 port map( A => n2739, B => n8110, C => n2738, D => n8109, Z => 
                           n554);
   U4263 : AO4 port map( A => n2747, B => n8102, C => n2746, D => n8101, Z => 
                           n558);
   U4264 : AO4 port map( A => n2691, B => n8094, C => n2690, D => n8093, Z => 
                           n566);
   U4265 : AO4 port map( A => n2699, B => n8086, C => n2698, D => n8085, Z => 
                           n570);
   U4266 : AO4 port map( A => n2707, B => n8078, C => n2706, D => n8077, Z => 
                           n574);
   U4267 : AO4 port map( A => n2715, B => n8070, C => n2714, D => n8069, Z => 
                           n578);
   U4268 : AO4 port map( A => n2788, B => n8126, C => n2787, D => n8125, Z => 
                           n590);
   U4269 : AO4 port map( A => n2796, B => n8118, C => n2795, D => n8117, Z => 
                           n594);
   U4270 : AO4 port map( A => n2804, B => n8110, C => n2803, D => n8109, Z => 
                           n598);
   U4271 : AO4 port map( A => n2812, B => n8102, C => n2811, D => n8101, Z => 
                           n602);
   U4272 : AO4 port map( A => n2756, B => n8094, C => n2755, D => n8093, Z => 
                           n610);
   U4273 : AO4 port map( A => n2764, B => n8086, C => n2763, D => n8085, Z => 
                           n614);
   U4274 : AO4 port map( A => n2772, B => n8078, C => n2771, D => n8077, Z => 
                           n618);
   U4275 : AO4 port map( A => n2780, B => n8070, C => n2779, D => n8069, Z => 
                           n622);
   U4276 : AO4 port map( A => n2852, B => n8126, C => n2851, D => n8125, Z => 
                           n634);
   U4277 : AO4 port map( A => n2860, B => n8118, C => n2859, D => n8117, Z => 
                           n638);
   U4278 : AO4 port map( A => n2868, B => n8110, C => n2867, D => n8109, Z => 
                           n642);
   U4279 : AO4 port map( A => n2876, B => n8102, C => n2875, D => n8101, Z => 
                           n646);
   U4280 : AO4 port map( A => n2820, B => n8094, C => n2819, D => n8093, Z => 
                           n654);
   U4281 : AO4 port map( A => n2828, B => n8086, C => n2827, D => n8085, Z => 
                           n658);
   U4282 : AO4 port map( A => n2836, B => n8078, C => n2835, D => n8077, Z => 
                           n662);
   U4283 : AO4 port map( A => n2844, B => n8070, C => n2843, D => n8069, Z => 
                           n666);
   U4284 : AO4 port map( A => n2916, B => n8126, C => n2915, D => n8125, Z => 
                           n678);
   U4285 : AO4 port map( A => n2924, B => n8118, C => n2923, D => n8117, Z => 
                           n682);
   U4286 : AO4 port map( A => n2932, B => n8110, C => n2931, D => n8109, Z => 
                           n686);
   U4287 : AO4 port map( A => n2940, B => n8102, C => n2939, D => n8101, Z => 
                           n690);
   U4288 : AO4 port map( A => n2884, B => n8094, C => n2883, D => n8093, Z => 
                           n698);
   U4289 : AO4 port map( A => n2892, B => n8086, C => n2891, D => n8085, Z => 
                           n702);
   U4290 : AO4 port map( A => n2900, B => n8078, C => n2899, D => n8077, Z => 
                           n706);
   U4291 : AO4 port map( A => n2908, B => n8070, C => n2907, D => n8069, Z => 
                           n710);
   U4292 : AO4 port map( A => n2980, B => n8126, C => n2979, D => n8125, Z => 
                           n721);
   U4293 : AO4 port map( A => n2988, B => n8118, C => n2987, D => n8117, Z => 
                           n725);
   U4294 : AO4 port map( A => n2996, B => n8110, C => n2995, D => n8109, Z => 
                           n729);
   U4295 : AO4 port map( A => n3004, B => n8102, C => n3003, D => n8101, Z => 
                           n733);
   U4296 : AO4 port map( A => n2948, B => n8094, C => n2947, D => n8093, Z => 
                           n741);
   U4297 : AO4 port map( A => n2956, B => n8086, C => n2955, D => n8085, Z => 
                           n745);
   U4298 : AO4 port map( A => n2964, B => n8078, C => n2963, D => n8077, Z => 
                           n749);
   U4299 : AO4 port map( A => n2972, B => n8070, C => n2971, D => n8069, Z => 
                           n753);
   U4300 : AO4 port map( A => n3044, B => n8126, C => n3043, D => n8125, Z => 
                           n765);
   U4301 : AO4 port map( A => n3052, B => n8118, C => n3051, D => n8117, Z => 
                           n769);
   U4302 : AO4 port map( A => n3060, B => n8110, C => n3059, D => n8109, Z => 
                           n773);
   U4303 : AO4 port map( A => n3068, B => n8102, C => n3067, D => n8101, Z => 
                           n777);
   U4304 : AO4 port map( A => n3012, B => n8094, C => n3011, D => n8093, Z => 
                           n785);
   U4305 : AO4 port map( A => n3020, B => n8086, C => n3019, D => n8085, Z => 
                           n789);
   U4306 : AO4 port map( A => n3028, B => n8078, C => n3027, D => n8077, Z => 
                           n793);
   U4307 : AO4 port map( A => n3036, B => n8070, C => n3035, D => n8069, Z => 
                           n797);
   U4308 : AO4 port map( A => n3108, B => n8126, C => n3107, D => n8125, Z => 
                           n809);
   U4309 : AO4 port map( A => n3116, B => n8118, C => n3115, D => n8117, Z => 
                           n813);
   U4310 : AO4 port map( A => n3124, B => n8110, C => n3123, D => n8109, Z => 
                           n817);
   U4311 : AO4 port map( A => n3132, B => n8102, C => n3131, D => n8101, Z => 
                           n821);
   U4312 : AO4 port map( A => n3076, B => n8094, C => n3075, D => n8093, Z => 
                           n829);
   U4313 : AO4 port map( A => n3084, B => n8086, C => n3083, D => n8085, Z => 
                           n833);
   U4314 : AO4 port map( A => n3092, B => n8078, C => n3091, D => n8077, Z => 
                           n837);
   U4315 : AO4 port map( A => n3100, B => n8070, C => n3099, D => n8069, Z => 
                           n841);
   U4316 : AO4 port map( A => n3172, B => n8126, C => n3171, D => n8125, Z => 
                           n853);
   U4317 : AO4 port map( A => n3180, B => n8118, C => n3179, D => n8117, Z => 
                           n857);
   U4318 : AO4 port map( A => n3188, B => n8110, C => n3187, D => n8109, Z => 
                           n861);
   U4319 : AO4 port map( A => n3196, B => n8102, C => n3195, D => n8101, Z => 
                           n865);
   U4320 : AO4 port map( A => n3140, B => n8094, C => n3139, D => n8093, Z => 
                           n873);
   U4321 : AO4 port map( A => n3148, B => n8086, C => n3147, D => n8085, Z => 
                           n877);
   U4322 : AO4 port map( A => n3156, B => n8078, C => n3155, D => n8077, Z => 
                           n881);
   U4323 : AO4 port map( A => n3164, B => n8070, C => n3163, D => n8069, Z => 
                           n885);
   U4324 : AO4 port map( A => n3236, B => n8126, C => n3235, D => n8125, Z => 
                           n896);
   U4325 : AO4 port map( A => n3244, B => n8118, C => n3243, D => n8117, Z => 
                           n900);
   U4326 : AO4 port map( A => n3252, B => n8110, C => n3251, D => n8109, Z => 
                           n904);
   U4327 : AO4 port map( A => n3260, B => n8102, C => n3259, D => n8101, Z => 
                           n908);
   U4328 : AO4 port map( A => n3204, B => n8094, C => n3203, D => n8093, Z => 
                           n916);
   U4329 : AO4 port map( A => n3212, B => n8086, C => n3211, D => n8085, Z => 
                           n920);
   U4330 : AO4 port map( A => n3220, B => n8078, C => n3219, D => n8077, Z => 
                           n924);
   U4331 : AO4 port map( A => n3228, B => n8070, C => n3227, D => n8069, Z => 
                           n928);
   U4332 : AO4 port map( A => n3300, B => n8126, C => n3299, D => n8125, Z => 
                           n940);
   U4333 : AO4 port map( A => n3308, B => n8118, C => n3307, D => n8117, Z => 
                           n944);
   U4334 : AO4 port map( A => n3316, B => n8110, C => n3315, D => n8109, Z => 
                           n948);
   U4335 : AO4 port map( A => n3324, B => n8102, C => n3323, D => n8101, Z => 
                           n952);
   U4336 : AO4 port map( A => n3268, B => n8094, C => n3267, D => n8093, Z => 
                           n960);
   U4337 : AO4 port map( A => n3276, B => n8086, C => n3275, D => n8085, Z => 
                           n964);
   U4338 : AO4 port map( A => n3284, B => n8078, C => n3283, D => n8077, Z => 
                           n968);
   U4339 : AO4 port map( A => n3292, B => n8070, C => n3291, D => n8069, Z => 
                           n972);
   U4340 : AO4 port map( A => n3364, B => n8126, C => n3363, D => n8125, Z => 
                           n984);
   U4341 : AO4 port map( A => n3372, B => n8118, C => n3371, D => n8117, Z => 
                           n988);
   U4342 : AO4 port map( A => n3380, B => n8110, C => n3379, D => n8109, Z => 
                           n992);
   U4343 : AO4 port map( A => n3388, B => n8102, C => n3387, D => n8101, Z => 
                           n996);
   U4344 : AO4 port map( A => n3332, B => n8094, C => n3331, D => n8093, Z => 
                           n1004);
   U4345 : AO4 port map( A => n3340, B => n8086, C => n3339, D => n8085, Z => 
                           n1008);
   U4346 : AO4 port map( A => n3348, B => n8078, C => n3347, D => n8077, Z => 
                           n1012);
   U4347 : AO4 port map( A => n3356, B => n8070, C => n3355, D => n8069, Z => 
                           n1016);
   U4348 : AO4 port map( A => n3428, B => n8126, C => n3427, D => n8125, Z => 
                           n1028);
   U4349 : AO4 port map( A => n3436, B => n8118, C => n3435, D => n8117, Z => 
                           n1032);
   U4350 : AO4 port map( A => n3444, B => n8110, C => n3443, D => n8109, Z => 
                           n1036);
   U4351 : AO4 port map( A => n3452, B => n8102, C => n3451, D => n8101, Z => 
                           n1040);
   U4352 : AO4 port map( A => n3396, B => n8094, C => n3395, D => n8093, Z => 
                           n1048);
   U4353 : AO4 port map( A => n3404, B => n8086, C => n3403, D => n8085, Z => 
                           n1052);
   U4354 : AO4 port map( A => n3412, B => n8078, C => n3411, D => n8077, Z => 
                           n1056);
   U4355 : AO4 port map( A => n3420, B => n8070, C => n3419, D => n8069, Z => 
                           n1060);
   U4356 : AO4 port map( A => n3492, B => n8126, C => n3491, D => n8125, Z => 
                           n1071);
   U4357 : AO4 port map( A => n3500, B => n8118, C => n3499, D => n8117, Z => 
                           n1075);
   U4358 : AO4 port map( A => n3508, B => n8110, C => n3507, D => n8109, Z => 
                           n1079);
   U4359 : AO4 port map( A => n3516, B => n8102, C => n3515, D => n8101, Z => 
                           n1083);
   U4360 : AO4 port map( A => n3460, B => n8094, C => n3459, D => n8093, Z => 
                           n1091);
   U4361 : AO4 port map( A => n3468, B => n8086, C => n3467, D => n8085, Z => 
                           n1095);
   U4362 : AO4 port map( A => n3476, B => n8078, C => n3475, D => n8077, Z => 
                           n1099);
   U4363 : AO4 port map( A => n3484, B => n8070, C => n3483, D => n8069, Z => 
                           n1103);
   U4364 : AO4 port map( A => n3556, B => n8126, C => n3555, D => n8125, Z => 
                           n1115);
   U4365 : AO4 port map( A => n3564, B => n8118, C => n3563, D => n8117, Z => 
                           n1119);
   U4366 : AO4 port map( A => n3572, B => n8110, C => n3571, D => n8109, Z => 
                           n1123);
   U4367 : AO4 port map( A => n3580, B => n8102, C => n3579, D => n8101, Z => 
                           n1127);
   U4368 : AO4 port map( A => n3524, B => n8094, C => n3523, D => n8093, Z => 
                           n1135);
   U4369 : AO4 port map( A => n3532, B => n8086, C => n3531, D => n8085, Z => 
                           n1139);
   U4370 : AO4 port map( A => n3540, B => n8078, C => n3539, D => n8077, Z => 
                           n1143);
   U4371 : AO4 port map( A => n3548, B => n8070, C => n3547, D => n8069, Z => 
                           n1147);
   U4372 : AO4 port map( A => n3620, B => n8126, C => n3619, D => n8125, Z => 
                           n1159);
   U4373 : AO4 port map( A => n3628, B => n8118, C => n3627, D => n8117, Z => 
                           n1163);
   U4374 : AO4 port map( A => n3636, B => n8110, C => n3635, D => n8109, Z => 
                           n1167);
   U4375 : AO4 port map( A => n3644, B => n8102, C => n3643, D => n8101, Z => 
                           n1171);
   U4376 : AO4 port map( A => n3588, B => n8094, C => n3587, D => n8093, Z => 
                           n1179);
   U4377 : AO4 port map( A => n3596, B => n8086, C => n3595, D => n8085, Z => 
                           n1183);
   U4378 : AO4 port map( A => n3604, B => n8078, C => n3603, D => n8077, Z => 
                           n1187);
   U4379 : AO4 port map( A => n3612, B => n8070, C => n3611, D => n8069, Z => 
                           n1191);
   U4380 : AO4 port map( A => n3684, B => n8126, C => n3683, D => n8125, Z => 
                           n1203);
   U4381 : AO4 port map( A => n3692, B => n8118, C => n3691, D => n8117, Z => 
                           n1207);
   U4382 : AO4 port map( A => n3700, B => n8110, C => n3699, D => n8109, Z => 
                           n1211);
   U4383 : AO4 port map( A => n3708, B => n8102, C => n3707, D => n8101, Z => 
                           n1215);
   U4384 : AO4 port map( A => n3652, B => n8094, C => n3651, D => n8093, Z => 
                           n1223);
   U4385 : AO4 port map( A => n3660, B => n8086, C => n3659, D => n8085, Z => 
                           n1227);
   U4386 : AO4 port map( A => n3668, B => n8078, C => n3667, D => n8077, Z => 
                           n1231);
   U4387 : AO4 port map( A => n3676, B => n8070, C => n3675, D => n8069, Z => 
                           n1235);
   U4388 : AO4 port map( A => n3748, B => n8126, C => n3747, D => n8125, Z => 
                           n1246);
   U4389 : AO4 port map( A => n3756, B => n8118, C => n3755, D => n8117, Z => 
                           n1250);
   U4390 : AO4 port map( A => n3764, B => n8110, C => n3763, D => n8109, Z => 
                           n1254);
   U4391 : AO4 port map( A => n3772, B => n8102, C => n3771, D => n8101, Z => 
                           n1258);
   U4392 : AO4 port map( A => n3716, B => n8094, C => n3715, D => n8093, Z => 
                           n1266);
   U4393 : AO4 port map( A => n3724, B => n8086, C => n3723, D => n8085, Z => 
                           n1270);
   U4394 : AO4 port map( A => n3732, B => n8078, C => n3731, D => n8077, Z => 
                           n1274);
   U4395 : AO4 port map( A => n3740, B => n8070, C => n3739, D => n8069, Z => 
                           n1278);
   U4396 : AO4 port map( A => n3812, B => n8126, C => n3811, D => n8125, Z => 
                           n1290);
   U4397 : AO4 port map( A => n3820, B => n8118, C => n3819, D => n8117, Z => 
                           n1294);
   U4398 : AO4 port map( A => n3828, B => n8110, C => n3827, D => n8109, Z => 
                           n1298);
   U4399 : AO4 port map( A => n3836, B => n8102, C => n3835, D => n8101, Z => 
                           n1302);
   U4400 : AO4 port map( A => n3780, B => n8094, C => n3779, D => n8093, Z => 
                           n1310);
   U4401 : AO4 port map( A => n3788, B => n8086, C => n3787, D => n8085, Z => 
                           n1314);
   U4402 : AO4 port map( A => n3796, B => n8078, C => n3795, D => n8077, Z => 
                           n1318);
   U4403 : AO4 port map( A => n3804, B => n8070, C => n3803, D => n8069, Z => 
                           n1322);
   U4404 : AO4 port map( A => n3876, B => n8126, C => n3875, D => n8125, Z => 
                           n1334);
   U4405 : AO4 port map( A => n3884, B => n8118, C => n3883, D => n8117, Z => 
                           n1338);
   U4406 : AO4 port map( A => n3892, B => n8110, C => n3891, D => n8109, Z => 
                           n1342);
   U4407 : AO4 port map( A => n3900, B => n8102, C => n3899, D => n8101, Z => 
                           n1346);
   U4408 : AO4 port map( A => n3844, B => n8094, C => n3843, D => n8093, Z => 
                           n1354);
   U4409 : AO4 port map( A => n3852, B => n8086, C => n3851, D => n8085, Z => 
                           n1358);
   U4410 : AO4 port map( A => n3860, B => n8078, C => n3859, D => n8077, Z => 
                           n1362);
   U4411 : AO4 port map( A => n3868, B => n8070, C => n3867, D => n8069, Z => 
                           n1366);
   U4412 : AO4 port map( A => n3940, B => n8126, C => n3939, D => n8125, Z => 
                           n1378);
   U4413 : AO4 port map( A => n3948, B => n8118, C => n3947, D => n8117, Z => 
                           n1382);
   U4414 : AO4 port map( A => n3956, B => n8110, C => n3955, D => n8109, Z => 
                           n1386);
   U4415 : AO4 port map( A => n3964, B => n8102, C => n3963, D => n8101, Z => 
                           n1390);
   U4416 : AO4 port map( A => n3908, B => n8094, C => n3907, D => n8093, Z => 
                           n1398);
   U4417 : AO4 port map( A => n3916, B => n8086, C => n3915, D => n8085, Z => 
                           n1402);
   U4418 : AO4 port map( A => n3924, B => n8078, C => n3923, D => n8077, Z => 
                           n1406);
   U4419 : AO4 port map( A => n3932, B => n8070, C => n3931, D => n8069, Z => 
                           n1410);
   U4420 : AO4 port map( A => n4004, B => n8126, C => n4003, D => n8125, Z => 
                           n1421);
   U4421 : AO4 port map( A => n4012, B => n8118, C => n4011, D => n8117, Z => 
                           n1425);
   U4422 : AO4 port map( A => n4020, B => n8110, C => n4019, D => n8109, Z => 
                           n1429);
   U4423 : AO4 port map( A => n4028, B => n8102, C => n4027, D => n8101, Z => 
                           n1433);
   U4424 : AO4 port map( A => n3972, B => n8094, C => n3971, D => n8093, Z => 
                           n1441);
   U4425 : AO4 port map( A => n3980, B => n8086, C => n3979, D => n8085, Z => 
                           n1445);
   U4426 : AO4 port map( A => n3988, B => n8078, C => n3987, D => n8077, Z => 
                           n1449);
   U4427 : AO4 port map( A => n3996, B => n8070, C => n3995, D => n8069, Z => 
                           n1453);
   U4428 : AO4 port map( A => n4068, B => n8126, C => n4067, D => n8125, Z => 
                           n1465);
   U4429 : AO4 port map( A => n4076, B => n8118, C => n4075, D => n8117, Z => 
                           n1469);
   U4430 : AO4 port map( A => n4084, B => n8110, C => n4083, D => n8109, Z => 
                           n1473);
   U4431 : AO4 port map( A => n4092, B => n8102, C => n4091, D => n8101, Z => 
                           n1477);
   U4432 : AO4 port map( A => n4036, B => n8094, C => n4035, D => n8093, Z => 
                           n1485);
   U4433 : AO4 port map( A => n4044, B => n8086, C => n4043, D => n8085, Z => 
                           n1489);
   U4434 : AO4 port map( A => n4052, B => n8078, C => n4051, D => n8077, Z => 
                           n1493);
   U4435 : AO4 port map( A => n4060, B => n8070, C => n4059, D => n8069, Z => 
                           n1497);
   U4436 : AO4 port map( A => n4132, B => n8126, C => n4131, D => n8125, Z => 
                           n1509);
   U4437 : AO4 port map( A => n4140, B => n8118, C => n4139, D => n8117, Z => 
                           n1513);
   U4438 : AO4 port map( A => n4148, B => n8110, C => n4147, D => n8109, Z => 
                           n1517);
   U4439 : AO4 port map( A => n4156, B => n8102, C => n4155, D => n8101, Z => 
                           n1521);
   U4440 : AO4 port map( A => n4100, B => n8094, C => n4099, D => n8093, Z => 
                           n1529);
   U4441 : AO4 port map( A => n4108, B => n8086, C => n4107, D => n8085, Z => 
                           n1533);
   U4442 : AO4 port map( A => n4116, B => n8078, C => n4115, D => n8077, Z => 
                           n1537);
   U4443 : AO4 port map( A => n4124, B => n8070, C => n4123, D => n8069, Z => 
                           n1541);
   U4444 : AO4 port map( A => n4196, B => n8126, C => n4195, D => n8125, Z => 
                           n1553);
   U4445 : AO4 port map( A => n4204, B => n8118, C => n4203, D => n8117, Z => 
                           n1557);
   U4446 : AO4 port map( A => n4212, B => n8110, C => n4211, D => n8109, Z => 
                           n1561);
   U4447 : AO4 port map( A => n4220, B => n8102, C => n4219, D => n8101, Z => 
                           n1565);
   U4448 : AO4 port map( A => n4164, B => n8094, C => n4163, D => n8093, Z => 
                           n1573);
   U4449 : AO4 port map( A => n4172, B => n8086, C => n4171, D => n8085, Z => 
                           n1577);
   U4450 : AO4 port map( A => n4180, B => n8078, C => n4179, D => n8077, Z => 
                           n1581);
   U4451 : AO4 port map( A => n4188, B => n8070, C => n4187, D => n8069, Z => 
                           n1585);
   U4452 : AO4 port map( A => n4260, B => n8126, C => n4259, D => n8125, Z => 
                           n1597);
   U4453 : AO4 port map( A => n4268, B => n8118, C => n4267, D => n8117, Z => 
                           n1601);
   U4454 : AO4 port map( A => n4276, B => n8110, C => n4275, D => n8109, Z => 
                           n1605);
   U4455 : AO4 port map( A => n4284, B => n8102, C => n4283, D => n8101, Z => 
                           n1609);
   U4456 : AO4 port map( A => n4228, B => n8094, C => n4227, D => n8093, Z => 
                           n1617);
   U4457 : AO4 port map( A => n4236, B => n8086, C => n4235, D => n8085, Z => 
                           n1621);
   U4458 : AO4 port map( A => n4244, B => n8078, C => n4243, D => n8077, Z => 
                           n1625);
   U4459 : AO4 port map( A => n4252, B => n8070, C => n4251, D => n8069, Z => 
                           n1629);
   U4460 : AO4 port map( A => n4325, B => n8126, C => n4324, D => n8125, Z => 
                           n1641);
   U4461 : AO4 port map( A => n4333, B => n8118, C => n4332, D => n8117, Z => 
                           n1645);
   U4462 : AO4 port map( A => n4341, B => n8110, C => n4340, D => n8109, Z => 
                           n1649);
   U4463 : AO4 port map( A => n4349, B => n8102, C => n4348, D => n8101, Z => 
                           n1653);
   U4464 : AO4 port map( A => n4293, B => n8094, C => n4292, D => n8093, Z => 
                           n1661);
   U4465 : AO4 port map( A => n4301, B => n8086, C => n4300, D => n8085, Z => 
                           n1665);
   U4466 : AO4 port map( A => n4309, B => n8078, C => n4308, D => n8077, Z => 
                           n1669);
   U4467 : AO4 port map( A => n4317, B => n8070, C => n4316, D => n8069, Z => 
                           n1673);
   U4468 : AO4 port map( A => n4389, B => n8126, C => n4388, D => n8125, Z => 
                           n1685);
   U4470 : AO4 port map( A => n4397, B => n8118, C => n4396, D => n8117, Z => 
                           n1689);
   U4471 : AO4 port map( A => n4405, B => n8110, C => n4404, D => n8109, Z => 
                           n1693);
   U4472 : AO4 port map( A => n4413, B => n8102, C => n4412, D => n8101, Z => 
                           n1697);
   U4473 : AO4 port map( A => n4357, B => n8094, C => n4356, D => n8093, Z => 
                           n1705);
   U4474 : AO4 port map( A => n4365, B => n8086, C => n4364, D => n8085, Z => 
                           n1709);
   U4475 : AO4 port map( A => n4373, B => n8078, C => n4372, D => n8077, Z => 
                           n1713);
   U4476 : AO4 port map( A => n4381, B => n8070, C => n4380, D => n8069, Z => 
                           n1717);
   U4477 : AO4 port map( A => n4453, B => n8126, C => n4452, D => n8125, Z => 
                           n1729);
   U4478 : AO4 port map( A => n4461, B => n8118, C => n4460, D => n8117, Z => 
                           n1733);
   U4479 : AO4 port map( A => n4469, B => n8110, C => n4468, D => n8109, Z => 
                           n1737);
   U4480 : AO4 port map( A => n4477, B => n8102, C => n4476, D => n8101, Z => 
                           n1741);
   U4481 : AO4 port map( A => n4421, B => n8094, C => n4420, D => n8093, Z => 
                           n1749_port);
   U4482 : AO4 port map( A => n4429, B => n8086, C => n4428, D => n8085, Z => 
                           n1753_port);
   U4483 : AO4 port map( A => n4437, B => n8078, C => n4436, D => n8077, Z => 
                           n1757);
   U4484 : AO4 port map( A => n4445, B => n8070, C => n4444, D => n8069, Z => 
                           n1761);
   U4485 : AO4 port map( A => n4517, B => n8126, C => n4516, D => n8125, Z => 
                           n1772);
   U4486 : AO4 port map( A => n4525, B => n8118, C => n4524, D => n8117, Z => 
                           n1785);
   U4487 : AO4 port map( A => n4533, B => n8110, C => n4532, D => n8109, Z => 
                           n1795);
   U4488 : AO4 port map( A => n4541, B => n8102, C => n4540, D => n8101, Z => 
                           n1802);
   U4489 : AO4 port map( A => n4485, B => n8094, C => n4484, D => n8093, Z => 
                           n1814);
   U4490 : AO4 port map( A => n4493, B => n8086, C => n4492, D => n8085, Z => 
                           n1821);
   U4491 : AO4 port map( A => n4501, B => n8078, C => n4500, D => n8077, Z => 
                           n1827);
   U4492 : AO4 port map( A => n4509, B => n8070, C => n4508, D => n8069, Z => 
                           n1838);
   U4493 : AO4 port map( A => n6644, B => n260, C => n1919, D => n262, Z => 
                           n6703);
   U4495 : AO4 port map( A => n6645, B => n260, C => n1932, D => n262, Z => 
                           n6704);
   U4496 : AO4 port map( A => n6646, B => n260, C => n1947, D => n262, Z => 
                           n6705);
   U4497 : AO4 port map( A => n6647, B => n260, C => n1986, D => n262, Z => 
                           n6706);
   U4498 : EOI port map( A => n6648, B => i_INTERN_ADDR_RD0_0_port, Z => n2092)
                           ;
   U4499 : AO4 port map( A => n6649, B => n260, C => i_INTERN_ADDR_RD0_0_port, 
                           D => n262, Z => n6708);
   U4500 : AO7 port map( A => n6659, B => n8163, C => n8300, Z => n155);
   U4501 : EON1 port map( A => n317, B => n8301, C => N1751, D => n2482, Z => 
                           n6655);
   U4502 : EON1 port map( A => n375, B => n8301, C => N1750, D => n2482, Z => 
                           n6654);
   U4503 : EON1 port map( A => n365, B => n8301, C => N1749, D => n2482, Z => 
                           n6653);
   U4504 : EOI port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => N1748);
   U4505 : EON1 port map( A => n1985, B => n8301, C => n1985, D => n2482, Z => 
                           n6651);
   U4506 : AO2 port map( A => n2483, B => v_CALCULATION_CNTR_7_port, C => N1754
                           , D => n2482, Z => n2486);
   U4507 : NR3 port map( A => n2462, B => n6640, C => i_SRAM_ADDR_WR0_4_port, Z
                           => n2464);
   U4508 : NR3 port map( A => n2462, B => n6639, C => i_SRAM_ADDR_WR0_3_port, Z
                           => n2465);
   U4509 : NR3 port map( A => i_SRAM_ADDR_WR0_0_port, B => n6641, C => 
                           i_SRAM_ADDR_WR0_1_port, Z => n2457);
   U4510 : NR3 port map( A => n6643, B => n6641, C => i_SRAM_ADDR_WR0_1_port, Z
                           => n2458);
   U4511 : NR3 port map( A => n6642, B => n6641, C => i_SRAM_ADDR_WR0_0_port, Z
                           => n2459);
   U4512 : AO2 port map( A => n177, B => n228, C => n8281, D => n229, Z => n227
                           );
   U4513 : AO2 port map( A => n177, B => n178, C => n8281, D => n179, Z => n176
                           );
   U4514 : ND3 port map( A => n363, B => n1918, C => n6663, Z => n180);
   U4515 : NR3 port map( A => n6640, B => n6639, C => n2462, Z => n2466);
   U4516 : ND2I port map( A => n6659, B => n8300, Z => n65);
   U4517 : EON1 port map( A => n8284, B => n289, C => n363, D => n287, Z => 
                           n6713);
   U4518 : AO4 port map( A => n6663, B => n8283, C => n290, D => n8284, Z => 
                           n6714);
   U4520 : EON1 port map( A => n8284, B => n291, C => n1921, D => n292, Z => 
                           n6715);
   U4521 : AO7 port map( A => n65, B => n280, C => n8283, Z => n292);
   U4522 : NR3 port map( A => n6641, B => n6642, C => n6643, Z => n2460);
   U4523 : AO6 port map( A => n2488, B => n2487, C => n336, Z => n315);
   U4524 : AO6 port map( A => n8299, B => n4548, C => RESET_I, Z => n246);
   U4525 : AO4 port map( A => n6659, B => n281, C => n8215, D => n282, Z => 
                           n6711);
   U4526 : AO7 port map( A => n8287, B => n1921, C => n8142, Z => n284);
   U4527 : AO6 port map( A => n1921, B => n6663, C => n207, Z => n205);
   U4528 : AO7 port map( A => n2491, B => n8301, C => n249, Z => n6702);
   U4529 : AO3 port map( A => n157, B => n250, C => n8300, D => n8140, Z => 
                           n249);
   U4530 : AO4 port map( A => n2489, B => n272, C => n8216, D => n277, Z => 
                           n6710);
   U4531 : ND3 port map( A => n280, B => n8142, C => n6660, Z => n279);
   U4532 : AO2 port map( A => KEY_I(0), B => n8189, C => n328, D => 
                           v_KEY32_IN_24_port, Z => n326);
   U4533 : AO2 port map( A => KEY_I(1), B => n8189, C => n328, D => 
                           v_KEY32_IN_25_port, Z => n329);
   U4534 : AO2 port map( A => KEY_I(2), B => n8189, C => n328, D => 
                           v_KEY32_IN_26_port, Z => n330);
   U4535 : AO2 port map( A => KEY_I(3), B => n8189, C => n328, D => 
                           v_KEY32_IN_27_port, Z => n331);
   U4536 : AO2 port map( A => KEY_I(4), B => n8189, C => n328, D => 
                           v_KEY32_IN_28_port, Z => n332);
   U4537 : AO2 port map( A => KEY_I(5), B => n8189, C => n328, D => 
                           v_KEY32_IN_29_port, Z => n333);
   U4538 : AO2 port map( A => KEY_I(6), B => n8189, C => n328, D => 
                           v_KEY32_IN_30_port, Z => n334);
   U4539 : AO2 port map( A => KEY_I(7), B => n8189, C => n328, D => 
                           v_KEY32_IN_31_port, Z => n335);
   U4540 : AN3 port map( A => n8299, B => n2488, C => n2487, Z => n296);
   U4541 : AO2 port map( A => n6663, B => n215, C => n6660, D => n290, Z => 
                           n214);
   U4542 : AO4 port map( A => n6638, B => n237, C => n1920, D => n239, Z => 
                           n6701);
   U4543 : AO2 port map( A => n2298, B => KEY_I(0), C => n1909, D => 
                           v_KEY32_IN_0_port, Z => n295);
   U4545 : AO2 port map( A => n2298, B => KEY_I(1), C => n1909, D => 
                           v_KEY32_IN_1_port, Z => n298);
   U4546 : AO2 port map( A => n2298, B => KEY_I(2), C => n1909, D => 
                           v_KEY32_IN_2_port, Z => n299);
   U4547 : AO2 port map( A => n2298, B => KEY_I(3), C => n1909, D => 
                           v_KEY32_IN_3_port, Z => n300);
   U4549 : AO2 port map( A => n2298, B => KEY_I(4), C => n1909, D => 
                           v_KEY32_IN_4_port, Z => n301);
   U4550 : AO2 port map( A => n296, B => KEY_I(5), C => n1909, D => 
                           v_KEY32_IN_5_port, Z => n302);
   U4551 : AO2 port map( A => n296, B => KEY_I(6), C => n1909, D => 
                           v_KEY32_IN_6_port, Z => n303);
   U4553 : AO2 port map( A => n296, B => KEY_I(7), C => n1909, D => 
                           v_KEY32_IN_7_port, Z => n304);
   U4554 : AO2 port map( A => KEY_I(0), B => n1910, C => n2296, D => 
                           v_KEY32_IN_8_port, Z => n305);
   U4555 : AO2 port map( A => KEY_I(1), B => n1910, C => n2296, D => 
                           v_KEY32_IN_9_port, Z => n308);
   U4557 : AO2 port map( A => KEY_I(2), B => n1910, C => n2296, D => 
                           v_KEY32_IN_10_port, Z => n309);
   U4558 : AO2 port map( A => KEY_I(3), B => n1910, C => n2296, D => 
                           v_KEY32_IN_11_port, Z => n310);
   U4559 : AO2 port map( A => KEY_I(4), B => n1910, C => n2296, D => 
                           v_KEY32_IN_12_port, Z => n311);
   U4561 : AO2 port map( A => KEY_I(5), B => n1910, C => n2296, D => 
                           v_KEY32_IN_13_port, Z => n312);
   U4562 : AO2 port map( A => KEY_I(6), B => n1910, C => n2296, D => 
                           v_KEY32_IN_14_port, Z => n313);
   U4563 : AO2 port map( A => KEY_I(7), B => n1910, C => n2296, D => 
                           v_KEY32_IN_15_port, Z => n314);
   U4564 : AO2 port map( A => KEY_I(0), B => n8206, C => n318, D => 
                           v_KEY32_IN_16_port, Z => n316);
   U4565 : AO2 port map( A => KEY_I(1), B => n8206, C => n318, D => 
                           v_KEY32_IN_17_port, Z => n319);
   U4566 : AO2 port map( A => KEY_I(2), B => n8206, C => n318, D => 
                           v_KEY32_IN_18_port, Z => n320);
   U4567 : AO2 port map( A => KEY_I(3), B => n8206, C => n318, D => 
                           v_KEY32_IN_19_port, Z => n321);
   U4568 : AO2 port map( A => KEY_I(4), B => n8206, C => n318, D => 
                           v_KEY32_IN_20_port, Z => n322);
   U4569 : AO2 port map( A => KEY_I(5), B => n8206, C => n318, D => 
                           v_KEY32_IN_21_port, Z => n323);
   U4570 : AO2 port map( A => KEY_I(6), B => n8206, C => n318, D => 
                           v_KEY32_IN_22_port, Z => n324);
   U4571 : AO2 port map( A => KEY_I(7), B => n8206, C => n318, D => 
                           v_KEY32_IN_23_port, Z => n325);
   U4572 : AO6 port map( A => n8142, B => n283, C => RESET_I, Z => n278);
   U4573 : AO7 port map( A => n290, B => n190, C => n6660, Z => n197);
   U4574 : AO4 port map( A => n6639, B => n237, C => n1943, D => n239, Z => 
                           n6696);
   U4575 : AO4 port map( A => n6640, B => n237, C => n1953, D => n239, Z => 
                           n6697);
   U4576 : AO4 port map( A => n6641, B => n237, C => n1989, D => n239, Z => 
                           n6698);
   U4577 : EOI port map( A => n6642, B => i_SRAM_ADDR_WR0_0_port, Z => n2095);
   U4579 : AO4 port map( A => n6643, B => n237, C => i_SRAM_ADDR_WR0_0_port, D 
                           => n239, Z => n6700);
   U4584 : AO6 port map( A => VALID_KEY_I, B => n4548, C => RESET_I, Z => n245)
                           ;
   U4587 : AO6 port map( A => n190, B => n6660, C => n6663, Z => n189);
   U4588 : AO4 port map( A => n2487, B => n8142, C => n336, D => n288, Z => 
                           n6749);
   U4589 : AO4 port map( A => n2488, B => n337, C => n358, D => n338, Z => 
                           n6748);
   U4590 : AO6 port map( A => n2487, B => VALID_KEY_I, C => n8161, Z => n337);
   U4591 : AO7 port map( A => n4548, B => n8140, C => n336, Z => n4589);
   U4592 : IVDA port map( A => n236, Y => n_3136, Z => n2111);
   U4593 : IVI port map( A => n1888, Z => n8257);
   U4596 : AO4 port map( A => n8257, B => n2279, C => n2065, D => n2262, Z => 
                           n2063);
   U4598 : AO2 port map( A => v_TEMP_VECTOR_8_port, B => n364, C => 
                           v_TEMP_VECTOR_0_port, D => n2247, Z => n2264);
   U4599 : NR3 port map( A => n364, B => n156, C => n157, Z => n232);
   U4600 : AO2 port map( A => v_TEMP_VECTOR_14_port, B => n364, C => 
                           v_TEMP_VECTOR_6_port, D => n2247, Z => n2245);
   U4601 : AO2 port map( A => v_TEMP_VECTOR_13_port, B => n364, C => 
                           v_TEMP_VECTOR_5_port, D => n2247, Z => n2266);
   U4602 : AO2 port map( A => v_TEMP_VECTOR_9_port, B => n364, C => 
                           v_TEMP_VECTOR_1_port, D => n2247, Z => n2272);
   U4603 : ND3 port map( A => n2082, B => n2147, C => n2040, Z => n2146);
   U4604 : IVI port map( A => n2077, Z => n8251);
   U4605 : AO3 port map( A => n1884, B => n1869, C => n1945, D => n1946, Z => 
                           n1944);
   U4606 : AO4 port map( A => n8242, B => n2288, C => n2053, D => n1869, Z => 
                           n2052);
   U4607 : AO6 port map( A => n8260, B => n1916, C => n2185, Z => n2176);
   U4608 : AO2 port map( A => n1860, B => n8260, C => n2114, D => n378, Z => 
                           n2165);
   U4609 : AO1 port map( A => n8260, B => n2127, C => n2203, D => n2204, Z => 
                           n2195);
   U4610 : AO2 port map( A => n2128, B => n368, C => n8260, D => n2065, Z => 
                           n2220);
   U4611 : AO2 port map( A => n8260, B => n2010, C => n2005, D => n2011, Z => 
                           n1998);
   U4612 : EO1 port map( A => n2005, B => n2082, C => n2083, D => n1869, Z => 
                           n2070);
   U4613 : AO7 port map( A => n1923, B => n2162, C => n1869, Z => n2253);
   U4614 : AO6 port map( A => n1869, B => n2161, C => n8250, Z => n2160);
   U4615 : AO2 port map( A => n8224, B => n8262, C => n8230, D => n8260, Z => 
                           n2034);
   U4616 : AO2 port map( A => n1895, B => n2035, C => n8267, D => n1898, Z => 
                           n1893);
   U4617 : AO1 port map( A => n8250, B => n2035, C => n2231, D => n1990, Z => 
                           n2230);
   U4618 : IVDA port map( A => n1935, Y => n370, Z => n2189);
   U4619 : AO3 port map( A => n8252, B => n2290, C => n1941, D => n2150, Z => 
                           n2117);
   U4620 : EON1 port map( A => n1863, B => n1957, C => n8264, D => n1886, Z => 
                           n2051);
   U4621 : AO2 port map( A => n8252, B => n1984, C => n1937, D => n369, Z => 
                           n1981);
   U4622 : AO1 port map( A => n1951, B => n1952, C => n8252, D => n8229, Z => 
                           n1950);
   U4623 : AO2 port map( A => n8252, B => n267, C => n8265, D => n2169, Z => 
                           n2023);
   U4624 : IVI port map( A => n297, Z => n2136);
   U4625 : AN3 port map( A => n2046, B => n8251, C => n2028, Z => n2042);
   U4626 : AO4 port map( A => n2174, B => n2060, C => n8232, D => n2234, Z => 
                           n2091);
   U4629 : AO1 port map( A => n2076, B => n2174, C => n2235, D => n1983, Z => 
                           n2229);
   U4631 : AO4 port map( A => n377, B => n2174, C => n8251, D => n2189, Z => 
                           n2106);
   U4633 : ND3 port map( A => n2027, B => n1908, C => n276, Z => n1901);
   U4635 : AO3 port map( A => n8230, B => n8244, C => n2174, D => n274, Z => 
                           n1902);
   U4637 : AO3 port map( A => n8227, B => n8258, C => n2174, D => n273, Z => 
                           n1913);
   U4639 : EON1 port map( A => n2174, B => n1957, C => n8265, D => n1975, Z => 
                           n1970);
   U4641 : AO2 port map( A => n2120, B => n2121, C => n4546, D => n8144, Z => 
                           n2119);
   U4643 : AO3 port map( A => n1868, B => n2189, C => n8270, D => n2215, Z => 
                           n2208);
   U4645 : AO4 port map( A => n1868, B => n1869, C => n1870, D => n2279, Z => 
                           n1866);
   U4647 : AO3 port map( A => n1967, B => n2210, C => n2211, D => n2212, Z => 
                           n2209);
   U4649 : AO3 port map( A => n1967, B => n1980, C => n1981, D => n1982, Z => 
                           n1979);
   U4651 : AO3 port map( A => n1967, B => n2093, C => n2094, D => n8254, Z => 
                           n2090);
   U4653 : AO3 port map( A => n2242, B => n1967, C => n2233, D => n2243, Z => 
                           n2238);
   U4655 : AO3 port map( A => n1858, B => n1967, C => n2022, D => n2023, Z => 
                           n2021);
   U4657 : NR3 port map( A => n1967, B => n8257, C => n2062, Z => n2182);
   U4659 : AO4 port map( A => n1880, B => n2189, C => n1967, D => n1972, Z => 
                           n1971);
   U4661 : AO4 port map( A => n2305, B => n2111, C => n8298, D => n253, Z => 
                           n250);
   U4663 : AO7 port map( A => n8282, B => n2111, C => n257, Z => n270);
   U4665 : AO7 port map( A => n2305, B => n2111, C => n58, Z => n156);
   U4667 : AO7 port map( A => n2129, B => n2130, C => n8274, Z => n2118);
   U4669 : AO4 port map( A => n2140, B => n1960, C => n167, D => n168, Z => 
                           n165);
   U4671 : AO4 port map( A => n2140, B => n1964, C => n187, D => n168, Z => 
                           n186);
   U4673 : AO4 port map( A => n2140, B => n1974, C => n195, D => n168, Z => 
                           n194);
   U4675 : AO4 port map( A => n2140, B => n1976, C => n203, D => n168, Z => 
                           n202);
   U4677 : AO4 port map( A => n2140, B => n1978, C => n212, D => n168, Z => 
                           n211);
   U4679 : AO4 port map( A => n2140, B => n1955, C => n220, D => n168, Z => 
                           n219);
   U4681 : AO2 port map( A => n2053, B => n368, C => n8247, D => n8261, Z => 
                           n2152);
   U4683 : AO4 port map( A => n2140, B => n1959, C => n175, D => n176, Z => 
                           n174);
   U4685 : AO4 port map( A => n175, B => n227, C => n2140, D => n1954, Z => 
                           n226);
   U4687 : AO1 port map( A => n1880, B => n8261, C => n2198, D => n2199, Z => 
                           n2197);
   U4689 : AO2 port map( A => n368, B => n1853, C => n8261, D => n1884, Z => 
                           n1945);
   U4691 : AO6 port map( A => n1860, B => n2085, C => n2108, Z => n2098);
   U4692 : EO1 port map( A => n2032, B => n8260, C => n2256, D => n2149, Z => 
                           n2150);
   U4693 : AO2 port map( A => n368, B => n2173, C => n2085, D => n2287, Z => 
                           n2172);
   U4694 : AO6 port map( A => n2134, B => n1994, C => n2256, Z => n2133);
   U4695 : AO7 port map( A => n2256, B => n1922, C => n2241, Z => n2239);
   U4696 : AO2 port map( A => n1860, B => n2085, C => n378, D => n2210, Z => 
                           n2219);
   U4697 : AO2 port map( A => n2002, B => n2037, C => n2085, D => n2003, Z => 
                           n2001);
   U4698 : AO4 port map( A => n2256, B => n1857, C => n1858, D => n2288, Z => 
                           n1855);
   U4699 : AO4 port map( A => n1963, B => n2256, C => n1869, D => n1980, Z => 
                           n2126);
   U4700 : AO4 port map( A => n2287, B => n2256, C => n2262, D => n2088, Z => 
                           n2087);
   U4701 : EO1 port map( A => n1870, B => n8261, C => n2256, D => n2079, Z => 
                           n2157);
   U4702 : EO1 port map( A => n2085, B => n2083, C => n2262, D => n2109, Z => 
                           n2251);
   U4703 : AO4 port map( A => n8257, B => n2256, C => n8243, D => n2279, Z => 
                           n2073);
   U4704 : AO3 port map( A => n8230, B => n1931, C => n2151, D => n2152, Z => 
                           n2116);
   U4705 : AO4 port map( A => n2110, B => n1931, C => n2279, D => n2053, Z => 
                           n2167);
   U4706 : AO3 port map( A => n2032, B => n1931, C => n8248, D => n2034, Z => 
                           n2017);
   U4707 : AO4 port map( A => n2107, B => n1931, C => n1869, D => n2259, Z => 
                           n2258);
   U4708 : AO4 port map( A => n1931, B => n1922, C => n1863, D => n2186, Z => 
                           n2185);
   U4709 : AO4 port map( A => n1931, B => n1934, C => n2279, D => n2127, Z => 
                           n2203);
   U4710 : AO4 port map( A => n2008, B => n1863, C => n2147, D => n1931, Z => 
                           n2198);
   U4711 : AO3 port map( A => n1969, B => n2210, C => n2232, D => n2233, Z => 
                           n2231);
   U4712 : AO4 port map( A => n1969, B => n1980, C => n1868, D => n2234, Z => 
                           n2103);
   U4713 : AO3 port map( A => n1969, B => n2007, C => n2024, D => n2025, Z => 
                           n2020);
   U4714 : EON1 port map( A => n1969, B => n1882, C => n8263, D => n2107, Z => 
                           n2105);
   U4715 : AO4 port map( A => n1969, B => n2054, C => n2128, D => n2234, Z => 
                           n2181);
   U4716 : AO4 port map( A => n8251, B => n1931, C => n2288, D => n1956, Z => 
                           n1949);
   U4717 : AO4 port map( A => n1967, B => n2114, C => n2031, D => n1969, Z => 
                           n2113);
   U4718 : ND2I port map( A => n2268, B => n2269, Z => n1896);
   U4719 : ND2I port map( A => n2274, B => n2275, Z => n1888);
   U4720 : AO1 port map( A => n8249, B => n8265, C => n2190, D => n2206, Z => 
                           n2188);
   U4721 : AO2 port map( A => n2483, B => v_CALCULATION_CNTR_5_port, C => N1752
                           , D => n2482, Z => n2484);
   U4722 : AO3 port map( A => n2049, B => n2288, C => n2070, D => n2071, Z => 
                           n2069);
   U4723 : AO2 port map( A => n2049, B => n8269, C => n8262, D => n1922, Z => 
                           n2151);
   U4724 : AO4 port map( A => n2078, B => n2290, C => n2124, D => n2077, Z => 
                           n2123);
   U4725 : AO4 port map( A => n2144, B => n1869, C => n1888, D => n2262, Z => 
                           n2202);
   U4726 : AO2 port map( A => n8261, B => n1886, C => n378, D => n1888, Z => 
                           n1873);
   U4727 : AO4 port map( A => n2290, B => n2010, C => n1861, D => n2077, Z => 
                           n2240);
   U4728 : ND3 port map( A => n2082, B => n2077, C => n8265, Z => n2094);
   U4729 : AO4 port map( A => n2049, B => n2035, C => n8267, D => n1853, Z => 
                           n2047);
   U4730 : AO4 port map( A => n2049, B => n1967, C => n2183, D => n2104, Z => 
                           n2102);
   U4731 : AO4 port map( A => n2262, B => n1882, C => n1863, D => n2077, Z => 
                           n2159);
   U4732 : AO2 port map( A => n8263, B => n2049, C => n2213, D => n8265, Z => 
                           n2263);
   U4733 : AO6 port map( A => n2077, B => n2027, C => n2078, Z => n1899);
   U4734 : AO2 port map( A => n2483, B => v_CALCULATION_CNTR_6_port, C => N1753
                           , D => n2482, Z => n2485);
   U4735 : AO2 port map( A => n8236, B => n8262, C => n2028, D => n2005, Z => 
                           n2221);
   U4736 : AO7 port map( A => n2028, B => n8223, C => n2085, Z => n2044);
   U4737 : AO4 port map( A => n2183, B => n2136, C => n1868, D => n2234, Z => 
                           n2184);
   U4738 : AO2 port map( A => n267, B => n2136, C => n8265, D => n2011, Z => 
                           n2236);
   U4739 : AO7 port map( A => n1879, B => n2028, C => n8263, Z => n2024);
   U4740 : AO4 port map( A => n274, B => n376, C => n2200, D => n1888, Z => 
                           n1908);
   U4741 : ND3 port map( A => n2043, B => n375, C => v_CALCULATION_CNTR_4_port,
                           Z => n257);
   U4742 : IVI port map( A => n379, Z => n2306);
   U4743 : IVI port map( A => n2312, Z => n2311);
   U4744 : IVI port map( A => n2451, Z => n2312);
   U4745 : IVI port map( A => n2318, Z => n2317);
   U4746 : IVI port map( A => n2450, Z => n2318);
   U4747 : IVI port map( A => n2324, Z => n2323);
   U4748 : IVI port map( A => n2449, Z => n2324);
   U4749 : IVI port map( A => n2330, Z => n2329);
   U4750 : IVI port map( A => n2448, Z => n2330);
   U4751 : IVI port map( A => n2336, Z => n2335);
   U4752 : IVI port map( A => n2447, Z => n2336);
   U4753 : IVI port map( A => n2342, Z => n2341);
   U4754 : IVI port map( A => n2446, Z => n2342);
   U4755 : IVI port map( A => n2348, Z => n2347);
   U4756 : IVI port map( A => n2445, Z => n2348);
   U4757 : IVI port map( A => n2354, Z => n2353);
   U4758 : IVI port map( A => n2444, Z => n2354);
   U4759 : IVI port map( A => n2360, Z => n2359);
   U4760 : IVI port map( A => n2443, Z => n2360);
   U4761 : IVI port map( A => n2366, Z => n2365);
   U4762 : IVI port map( A => n2442, Z => n2366);
   U4763 : IVI port map( A => n2372, Z => n2371);
   U4764 : IVI port map( A => n2441, Z => n2372);
   U4765 : IVI port map( A => n2378, Z => n2377);
   U4766 : IVI port map( A => n2440, Z => n2378);
   U4767 : IVI port map( A => n2384, Z => n2383);
   U4768 : IVI port map( A => n2439, Z => n2384);
   U4769 : IVI port map( A => n2390, Z => n2389);
   U4770 : IVI port map( A => n2438, Z => n2390);
   U4771 : IVI port map( A => n2396, Z => n2395);
   U4772 : IVI port map( A => n2437, Z => n2396);
   U4773 : IVI port map( A => n2402, Z => n2401);
   U4774 : IVI port map( A => n2436, Z => n2402);
   U4775 : IVI port map( A => n2408, Z => n2407);
   U4776 : IVI port map( A => n2435, Z => n2408);
   U4777 : IVI port map( A => n2414, Z => n2413);
   U4778 : IVI port map( A => n2434, Z => n2414);
   U4779 : IVI port map( A => n2420, Z => n2419);
   U4780 : IVI port map( A => n2433, Z => n2420);
   U4781 : IVI port map( A => n2481, Z => n2480);
   U4782 : IVI port map( A => n2432, Z => n2481);
   U4783 : IVI port map( A => n6657, Z => n6656);
   U4784 : IVI port map( A => n2431, Z => n6657);
   U4785 : IVI port map( A => n6720, Z => n6719);
   U4786 : IVI port map( A => n2430, Z => n6720);
   U4787 : IVI port map( A => n6726, Z => n6725);
   U4788 : IVI port map( A => n2429, Z => n6726);
   U4789 : IVI port map( A => n6732, Z => n6731);
   U4790 : IVI port map( A => n2428, Z => n6732);
   U4791 : IVI port map( A => n6738, Z => n6737);
   U4792 : IVI port map( A => n2427, Z => n6738);
   U4793 : IVI port map( A => n6744, Z => n6743);
   U4794 : IVI port map( A => n2426, Z => n6744);
   U4795 : IVI port map( A => n6752, Z => n6751);
   U4796 : IVI port map( A => n2425, Z => n6752);
   U4797 : IVI port map( A => n6758, Z => n6757);
   U4798 : IVI port map( A => n2424, Z => n6758);
   U4799 : IVI port map( A => n6764, Z => n6763);
   U4800 : IVI port map( A => n2423, Z => n6764);
   U4801 : IVI port map( A => n6770, Z => n6769);
   U4802 : IVI port map( A => n2422, Z => n6770);
   U4803 : IVI port map( A => n6776, Z => n6775);
   U4804 : IVI port map( A => n2421, Z => n6776);
   U4805 : IVI port map( A => n238, Z => n6777);
   U4806 : IVI port map( A => n238, Z => n6778);
   U4807 : IVI port map( A => n238, Z => n6779);
   U4808 : IVI port map( A => n238, Z => n6780);
   U4809 : IVI port map( A => n238, Z => n6781);
   U4810 : IVI port map( A => n238, Z => n6782);
   U4811 : IVI port map( A => n238, Z => n6783);
   U4812 : IVI port map( A => n238, Z => n6784);
   U4813 : IVI port map( A => n238, Z => n6785);
   U4814 : IVI port map( A => n238, Z => n6786);
   U4815 : IVI port map( A => n238, Z => n6787);
   U4816 : IVI port map( A => n238, Z => n6788);
   U4817 : IVI port map( A => n238, Z => n6789);
   U4818 : IVI port map( A => n238, Z => n6790);
   U4819 : IVI port map( A => n238, Z => n6791);
   U4820 : IVI port map( A => n238, Z => n6792);
   U4821 : IVI port map( A => n238, Z => n6793);
   U4822 : IVI port map( A => n6793, Z => n6796);
   U4823 : IVI port map( A => n235, Z => n6797);
   U4824 : IVI port map( A => n235, Z => n6798);
   U4825 : IVI port map( A => n235, Z => n6799);
   U4826 : IVI port map( A => n235, Z => n6800);
   U4827 : IVI port map( A => n235, Z => n6801);
   U4828 : IVI port map( A => n235, Z => n6802);
   U4829 : IVI port map( A => n235, Z => n6803);
   U4830 : IVI port map( A => n235, Z => n6804);
   U4831 : IVI port map( A => n235, Z => n6805);
   U4832 : IVI port map( A => n235, Z => n6806);
   U4833 : IVI port map( A => n235, Z => n6807);
   U4834 : IVI port map( A => n235, Z => n6808);
   U4835 : IVI port map( A => n235, Z => n6809);
   U4836 : IVI port map( A => n235, Z => n6810);
   U4837 : IVI port map( A => n235, Z => n6811);
   U4838 : IVI port map( A => n235, Z => n6812);
   U4839 : IVI port map( A => n235, Z => n6813);
   U4840 : IVI port map( A => n6813, Z => n6816);
   U4841 : IVI port map( A => n234, Z => n6817);
   U4842 : IVI port map( A => n234, Z => n6818);
   U4843 : IVI port map( A => n234, Z => n6819);
   U4844 : IVI port map( A => n234, Z => n6820);
   U4845 : IVI port map( A => n234, Z => n6821);
   U4846 : IVI port map( A => n234, Z => n6822);
   U4847 : IVI port map( A => n234, Z => n6823);
   U4848 : IVI port map( A => n234, Z => n6824);
   U4849 : IVI port map( A => n234, Z => n6825);
   U4850 : IVI port map( A => n234, Z => n6826);
   U4851 : IVI port map( A => n234, Z => n6827);
   U4852 : IVI port map( A => n234, Z => n6828);
   U4853 : IVI port map( A => n234, Z => n6829);
   U4854 : IVI port map( A => n234, Z => n6830);
   U4855 : IVI port map( A => n234, Z => n6831);
   U4856 : IVI port map( A => n234, Z => n6832);
   U4857 : IVI port map( A => n234, Z => n6833);
   U4858 : IVI port map( A => n6833, Z => n6836);
   U4859 : IVI port map( A => n233, Z => n6837);
   U4860 : IVI port map( A => n233, Z => n6838);
   U4861 : IVI port map( A => n233, Z => n6839);
   U4862 : IVI port map( A => n233, Z => n6840);
   U4863 : IVI port map( A => n233, Z => n6841);
   U4864 : IVI port map( A => n233, Z => n6842);
   U4865 : IVI port map( A => n233, Z => n6843);
   U4866 : IVI port map( A => n233, Z => n6844);
   U4867 : IVI port map( A => n233, Z => n6845);
   U4868 : IVI port map( A => n233, Z => n6846);
   U4869 : IVI port map( A => n233, Z => n6847);
   U4870 : IVI port map( A => n233, Z => n6848);
   U4871 : IVI port map( A => n233, Z => n6849);
   U4872 : IVI port map( A => n233, Z => n6850);
   U4873 : IVI port map( A => n233, Z => n6851);
   U4874 : IVI port map( A => n233, Z => n6852);
   U4875 : IVI port map( A => n233, Z => n6853);
   U4876 : IVI port map( A => n6853, Z => n6856);
   U4877 : IVI port map( A => n265, Z => n6857);
   U4878 : IVI port map( A => n265, Z => n6858);
   U4879 : IVI port map( A => n265, Z => n6859);
   U4880 : IVI port map( A => n265, Z => n6860);
   U4881 : IVI port map( A => n265, Z => n6861);
   U4882 : IVI port map( A => n265, Z => n6862);
   U4883 : IVI port map( A => n265, Z => n6863);
   U4884 : IVI port map( A => n265, Z => n6864);
   U4885 : IVI port map( A => n265, Z => n6865);
   U4886 : IVI port map( A => n265, Z => n6866);
   U4887 : IVI port map( A => n265, Z => n6867);
   U4888 : IVI port map( A => n265, Z => n6868);
   U4889 : IVI port map( A => n265, Z => n6869);
   U4890 : IVI port map( A => n265, Z => n6870);
   U4891 : IVI port map( A => n265, Z => n6871);
   U4892 : IVI port map( A => n265, Z => n6872);
   U4893 : IVI port map( A => n265, Z => n6873);
   U4894 : IVI port map( A => n6873, Z => n6876);
   U4895 : IVI port map( A => n264, Z => n6877);
   U4896 : IVI port map( A => n264, Z => n6878);
   U4897 : IVI port map( A => n264, Z => n6879);
   U4898 : IVI port map( A => n264, Z => n6880);
   U4899 : IVI port map( A => n264, Z => n6881);
   U4900 : IVI port map( A => n264, Z => n6882);
   U4901 : IVI port map( A => n264, Z => n6883);
   U4902 : IVI port map( A => n264, Z => n6884);
   U4903 : IVI port map( A => n264, Z => n6885);
   U4904 : IVI port map( A => n264, Z => n6886);
   U4905 : IVI port map( A => n264, Z => n6887);
   U4906 : IVI port map( A => n264, Z => n6888);
   U4907 : IVI port map( A => n264, Z => n6889);
   U4908 : IVI port map( A => n264, Z => n6890);
   U4909 : IVI port map( A => n264, Z => n6891);
   U4910 : IVI port map( A => n264, Z => n6892);
   U4911 : IVI port map( A => n264, Z => n6893);
   U4912 : IVI port map( A => n6893, Z => n6896);
   U4913 : IVI port map( A => n263, Z => n6897);
   U4914 : IVI port map( A => n263, Z => n6898);
   U4915 : IVI port map( A => n263, Z => n6899);
   U4916 : IVI port map( A => n263, Z => n6900);
   U4917 : IVI port map( A => n263, Z => n6901);
   U4918 : IVI port map( A => n263, Z => n6902);
   U4919 : IVI port map( A => n263, Z => n6903);
   U4920 : IVI port map( A => n263, Z => n6904);
   U4921 : IVI port map( A => n263, Z => n6905);
   U4922 : IVI port map( A => n263, Z => n6906);
   U4923 : IVI port map( A => n263, Z => n6907);
   U4924 : IVI port map( A => n263, Z => n6908);
   U4925 : IVI port map( A => n263, Z => n6909);
   U4926 : IVI port map( A => n263, Z => n6910);
   U4927 : IVI port map( A => n263, Z => n6911);
   U4928 : IVI port map( A => n263, Z => n6912);
   U4929 : IVI port map( A => n263, Z => n6913);
   U4930 : IVI port map( A => n6913, Z => n6916);
   U4931 : IVI port map( A => n261, Z => n6917);
   U4932 : IVI port map( A => n261, Z => n6918);
   U4933 : IVI port map( A => n261, Z => n6919);
   U4934 : IVI port map( A => n261, Z => n6920);
   U4935 : IVI port map( A => n261, Z => n6921);
   U4936 : IVI port map( A => n261, Z => n6922);
   U4937 : IVI port map( A => n261, Z => n6923);
   U4938 : IVI port map( A => n261, Z => n6924);
   U4939 : IVI port map( A => n261, Z => n6925);
   U4940 : IVI port map( A => n261, Z => n6926);
   U4941 : IVI port map( A => n261, Z => n6927);
   U4942 : IVI port map( A => n261, Z => n6928);
   U4943 : IVI port map( A => n261, Z => n6929);
   U4944 : IVI port map( A => n261, Z => n6930);
   U4945 : IVI port map( A => n261, Z => n6931);
   U4946 : IVI port map( A => n261, Z => n6932);
   U4947 : IVI port map( A => n261, Z => n6933);
   U4948 : IVI port map( A => n6933, Z => n6936);
   U4949 : IVI port map( A => n224, Z => n6937);
   U4950 : IVI port map( A => n224, Z => n6938);
   U4951 : IVI port map( A => n224, Z => n6939);
   U4952 : IVI port map( A => n224, Z => n6940);
   U4953 : IVI port map( A => n224, Z => n6941);
   U4954 : IVI port map( A => n224, Z => n6942);
   U4955 : IVI port map( A => n224, Z => n6943);
   U4956 : IVI port map( A => n224, Z => n6944);
   U4957 : IVI port map( A => n224, Z => n6945);
   U4958 : IVI port map( A => n224, Z => n6946);
   U4959 : IVI port map( A => n224, Z => n6947);
   U4960 : IVI port map( A => n224, Z => n6948);
   U4961 : IVI port map( A => n224, Z => n6949);
   U4962 : IVI port map( A => n224, Z => n6950);
   U4963 : IVI port map( A => n224, Z => n6951);
   U4964 : IVI port map( A => n224, Z => n6952);
   U4965 : IVI port map( A => n224, Z => n6953);
   U4966 : IVI port map( A => n6953, Z => n6956);
   U4967 : IVI port map( A => n221, Z => n6957);
   U4968 : IVI port map( A => n221, Z => n6958);
   U4969 : IVI port map( A => n221, Z => n6959);
   U4970 : IVI port map( A => n221, Z => n6960);
   U4971 : IVI port map( A => n221, Z => n6961);
   U4972 : IVI port map( A => n221, Z => n6962);
   U4973 : IVI port map( A => n221, Z => n6963);
   U4974 : IVI port map( A => n221, Z => n6964);
   U4975 : IVI port map( A => n221, Z => n6965);
   U4976 : IVI port map( A => n221, Z => n6966);
   U4977 : IVI port map( A => n221, Z => n6967);
   U4978 : IVI port map( A => n221, Z => n6968);
   U4979 : IVI port map( A => n221, Z => n6969);
   U4980 : IVI port map( A => n221, Z => n6970);
   U4981 : IVI port map( A => n221, Z => n6971);
   U4982 : IVI port map( A => n221, Z => n6972);
   U4983 : IVI port map( A => n221, Z => n6973);
   U4984 : IVI port map( A => n6973, Z => n6976);
   U4985 : IVI port map( A => n213, Z => n6977);
   U4986 : IVI port map( A => n213, Z => n6978);
   U4987 : IVI port map( A => n213, Z => n6979);
   U4988 : IVI port map( A => n213, Z => n6980);
   U4989 : IVI port map( A => n213, Z => n6981);
   U4990 : IVI port map( A => n213, Z => n6982);
   U4991 : IVI port map( A => n213, Z => n6983);
   U4992 : IVI port map( A => n213, Z => n6984);
   U4993 : IVI port map( A => n213, Z => n6985);
   U4994 : IVI port map( A => n213, Z => n6986);
   U4995 : IVI port map( A => n213, Z => n6987);
   U4996 : IVI port map( A => n213, Z => n6988);
   U4997 : IVI port map( A => n213, Z => n6989);
   U4998 : IVI port map( A => n213, Z => n6990);
   U4999 : IVI port map( A => n213, Z => n6991);
   U5000 : IVI port map( A => n213, Z => n6992);
   U5001 : IVI port map( A => n213, Z => n6993);
   U5002 : IVI port map( A => n6993, Z => n6996);
   U5003 : IVI port map( A => n206, Z => n6997);
   U5004 : IVI port map( A => n206, Z => n6998);
   U5005 : IVI port map( A => n206, Z => n6999);
   U5006 : IVI port map( A => n206, Z => n7000);
   U5007 : IVI port map( A => n206, Z => n7001);
   U5008 : IVI port map( A => n206, Z => n7002);
   U5009 : IVI port map( A => n206, Z => n7003);
   U5010 : IVI port map( A => n206, Z => n7004);
   U5011 : IVI port map( A => n206, Z => n7005);
   U5012 : IVI port map( A => n206, Z => n7006);
   U5013 : IVI port map( A => n206, Z => n7007);
   U5014 : IVI port map( A => n206, Z => n7008);
   U5015 : IVI port map( A => n206, Z => n7009);
   U5016 : IVI port map( A => n206, Z => n7010);
   U5017 : IVI port map( A => n206, Z => n7011);
   U5018 : IVI port map( A => n206, Z => n7012);
   U5019 : IVI port map( A => n206, Z => n7013);
   U5020 : IVI port map( A => n7013, Z => n7016);
   U5021 : IVI port map( A => n256, Z => n7017);
   U5022 : IVI port map( A => n256, Z => n7018);
   U5023 : IVI port map( A => n256, Z => n7019);
   U5024 : IVI port map( A => n256, Z => n7020);
   U5025 : IVI port map( A => n256, Z => n7021);
   U5026 : IVI port map( A => n256, Z => n7022);
   U5027 : IVI port map( A => n256, Z => n7023);
   U5028 : IVI port map( A => n256, Z => n7024);
   U5029 : IVI port map( A => n256, Z => n7025);
   U5030 : IVI port map( A => n256, Z => n7026);
   U5031 : IVI port map( A => n256, Z => n7027);
   U5032 : IVI port map( A => n256, Z => n7028);
   U5033 : IVI port map( A => n256, Z => n7029);
   U5034 : IVI port map( A => n256, Z => n7030);
   U5035 : IVI port map( A => n256, Z => n7031);
   U5036 : IVI port map( A => n256, Z => n7032);
   U5037 : IVI port map( A => n256, Z => n7033);
   U5038 : IVI port map( A => n7033, Z => n7036);
   U5039 : IVI port map( A => n255, Z => n7037);
   U5040 : IVI port map( A => n255, Z => n7038);
   U5041 : IVI port map( A => n255, Z => n7039);
   U5042 : IVI port map( A => n255, Z => n7040);
   U5043 : IVI port map( A => n255, Z => n7041);
   U5044 : IVI port map( A => n255, Z => n7042);
   U5045 : IVI port map( A => n255, Z => n7043);
   U5046 : IVI port map( A => n255, Z => n7044);
   U5047 : IVI port map( A => n255, Z => n7045);
   U5048 : IVI port map( A => n255, Z => n7046);
   U5049 : IVI port map( A => n255, Z => n7047);
   U5050 : IVI port map( A => n255, Z => n7048);
   U5051 : IVI port map( A => n255, Z => n7049);
   U5052 : IVI port map( A => n255, Z => n7050);
   U5053 : IVI port map( A => n255, Z => n7051);
   U5054 : IVI port map( A => n255, Z => n7052);
   U5055 : IVI port map( A => n255, Z => n7053);
   U5056 : IVI port map( A => n7053, Z => n7056);
   U5057 : IVI port map( A => n254, Z => n7057);
   U5058 : IVI port map( A => n254, Z => n7058);
   U5059 : IVI port map( A => n254, Z => n7059);
   U5060 : IVI port map( A => n254, Z => n7060);
   U5061 : IVI port map( A => n254, Z => n7061);
   U5062 : IVI port map( A => n254, Z => n7062);
   U5063 : IVI port map( A => n254, Z => n7063);
   U5064 : IVI port map( A => n254, Z => n7064);
   U5065 : IVI port map( A => n254, Z => n7065);
   U5066 : IVI port map( A => n254, Z => n7066);
   U5067 : IVI port map( A => n254, Z => n7067);
   U5068 : IVI port map( A => n254, Z => n7068);
   U5069 : IVI port map( A => n254, Z => n7069);
   U5070 : IVI port map( A => n254, Z => n7070);
   U5071 : IVI port map( A => n254, Z => n7071);
   U5072 : IVI port map( A => n254, Z => n7072);
   U5073 : IVI port map( A => n254, Z => n7073);
   U5074 : IVI port map( A => n7073, Z => n7076);
   U5075 : IVI port map( A => n252, Z => n7077);
   U5076 : IVI port map( A => n252, Z => n7078);
   U5077 : IVI port map( A => n252, Z => n7079);
   U5078 : IVI port map( A => n252, Z => n7080);
   U5079 : IVI port map( A => n252, Z => n7081);
   U5080 : IVI port map( A => n252, Z => n7082);
   U5081 : IVI port map( A => n252, Z => n7083);
   U5082 : IVI port map( A => n252, Z => n7084);
   U5083 : IVI port map( A => n252, Z => n7085);
   U5084 : IVI port map( A => n252, Z => n7086);
   U5085 : IVI port map( A => n252, Z => n7087);
   U5086 : IVI port map( A => n252, Z => n7088);
   U5087 : IVI port map( A => n252, Z => n7089);
   U5088 : IVI port map( A => n252, Z => n7090);
   U5089 : IVI port map( A => n252, Z => n7091);
   U5090 : IVI port map( A => n252, Z => n7092);
   U5091 : IVI port map( A => n252, Z => n7093);
   U5092 : IVI port map( A => n7093, Z => n7096);
   U5093 : IVI port map( A => n204, Z => n7097);
   U5094 : IVI port map( A => n204, Z => n7098);
   U5095 : IVI port map( A => n204, Z => n7099);
   U5096 : IVI port map( A => n204, Z => n7100);
   U5097 : IVI port map( A => n204, Z => n7101);
   U5098 : IVI port map( A => n204, Z => n7102);
   U5099 : IVI port map( A => n204, Z => n7103);
   U5100 : IVI port map( A => n204, Z => n7104);
   U5101 : IVI port map( A => n204, Z => n7105);
   U5102 : IVI port map( A => n204, Z => n7106);
   U5103 : IVI port map( A => n204, Z => n7107);
   U5104 : IVI port map( A => n204, Z => n7108);
   U5105 : IVI port map( A => n204, Z => n7109);
   U5106 : IVI port map( A => n204, Z => n7110);
   U5107 : IVI port map( A => n204, Z => n7111);
   U5108 : IVI port map( A => n204, Z => n7112);
   U5109 : IVI port map( A => n204, Z => n7113);
   U5110 : IVI port map( A => n7113, Z => n7116);
   U5111 : IVI port map( A => n198, Z => n7117);
   U5112 : IVI port map( A => n198, Z => n7118);
   U5113 : IVI port map( A => n198, Z => n7119);
   U5114 : IVI port map( A => n198, Z => n7120);
   U5115 : IVI port map( A => n198, Z => n7121);
   U5116 : IVI port map( A => n198, Z => n7122);
   U5117 : IVI port map( A => n198, Z => n7123);
   U5118 : IVI port map( A => n198, Z => n7124);
   U5119 : IVI port map( A => n198, Z => n7125);
   U5120 : IVI port map( A => n198, Z => n7126);
   U5121 : IVI port map( A => n198, Z => n7127);
   U5122 : IVI port map( A => n198, Z => n7128);
   U5123 : IVI port map( A => n198, Z => n7129);
   U5124 : IVI port map( A => n198, Z => n7130);
   U5125 : IVI port map( A => n198, Z => n7131);
   U5126 : IVI port map( A => n198, Z => n7132);
   U5127 : IVI port map( A => n198, Z => n7133);
   U5128 : IVI port map( A => n7133, Z => n7136);
   U5129 : IVI port map( A => n196, Z => n7137);
   U5130 : IVI port map( A => n196, Z => n7138);
   U5131 : IVI port map( A => n196, Z => n7139);
   U5132 : IVI port map( A => n196, Z => n7140);
   U5133 : IVI port map( A => n196, Z => n7141);
   U5134 : IVI port map( A => n196, Z => n7142);
   U5135 : IVI port map( A => n196, Z => n7143);
   U5136 : IVI port map( A => n196, Z => n7144);
   U5137 : IVI port map( A => n196, Z => n7145);
   U5138 : IVI port map( A => n196, Z => n7146);
   U5139 : IVI port map( A => n196, Z => n7147);
   U5140 : IVI port map( A => n196, Z => n7148);
   U5141 : IVI port map( A => n196, Z => n7149);
   U5142 : IVI port map( A => n196, Z => n7150);
   U5143 : IVI port map( A => n196, Z => n7151);
   U5144 : IVI port map( A => n196, Z => n7152);
   U5145 : IVI port map( A => n196, Z => n7153);
   U5146 : IVI port map( A => n7153, Z => n7156);
   U5147 : IVI port map( A => n188, Z => n7157);
   U5148 : IVI port map( A => n188, Z => n7158);
   U5149 : IVI port map( A => n188, Z => n7159);
   U5150 : IVI port map( A => n188, Z => n7160);
   U5151 : IVI port map( A => n188, Z => n7161);
   U5152 : IVI port map( A => n188, Z => n7162);
   U5153 : IVI port map( A => n188, Z => n7163);
   U5154 : IVI port map( A => n188, Z => n7164);
   U5155 : IVI port map( A => n188, Z => n7165);
   U5156 : IVI port map( A => n188, Z => n7166);
   U5157 : IVI port map( A => n188, Z => n7167);
   U5158 : IVI port map( A => n188, Z => n7168);
   U5159 : IVI port map( A => n188, Z => n7169);
   U5160 : IVI port map( A => n188, Z => n7170);
   U5161 : IVI port map( A => n188, Z => n7171);
   U5162 : IVI port map( A => n188, Z => n7172);
   U5163 : IVI port map( A => n188, Z => n7173);
   U5164 : IVI port map( A => n7173, Z => n7176);
   U5165 : IVI port map( A => n251, Z => n7177);
   U5166 : IVI port map( A => n251, Z => n7178);
   U5167 : IVI port map( A => n251, Z => n7179);
   U5168 : IVI port map( A => n251, Z => n7180);
   U5169 : IVI port map( A => n251, Z => n7181);
   U5170 : IVI port map( A => n251, Z => n7182);
   U5171 : IVI port map( A => n251, Z => n7183);
   U5172 : IVI port map( A => n251, Z => n7184);
   U5173 : IVI port map( A => n251, Z => n7185);
   U5174 : IVI port map( A => n251, Z => n7186);
   U5175 : IVI port map( A => n251, Z => n7187);
   U5176 : IVI port map( A => n251, Z => n7188);
   U5177 : IVI port map( A => n251, Z => n7189);
   U5178 : IVI port map( A => n251, Z => n7190);
   U5179 : IVI port map( A => n251, Z => n7191);
   U5180 : IVI port map( A => n251, Z => n7192);
   U5181 : IVI port map( A => n251, Z => n7193);
   U5182 : IVI port map( A => n7193, Z => n7196);
   U5183 : IVI port map( A => n248, Z => n7197);
   U5184 : IVI port map( A => n248, Z => n7198);
   U5185 : IVI port map( A => n248, Z => n7199);
   U5186 : IVI port map( A => n248, Z => n7200);
   U5187 : IVI port map( A => n248, Z => n7201);
   U5188 : IVI port map( A => n248, Z => n7202);
   U5189 : IVI port map( A => n248, Z => n7203);
   U5190 : IVI port map( A => n248, Z => n7204);
   U5191 : IVI port map( A => n248, Z => n7205);
   U5192 : IVI port map( A => n248, Z => n7206);
   U5193 : IVI port map( A => n248, Z => n7207);
   U5194 : IVI port map( A => n248, Z => n7208);
   U5195 : IVI port map( A => n248, Z => n7209);
   U5196 : IVI port map( A => n248, Z => n7210);
   U5197 : IVI port map( A => n248, Z => n7211);
   U5198 : IVI port map( A => n248, Z => n7212);
   U5199 : IVI port map( A => n248, Z => n7213);
   U5200 : IVI port map( A => n7213, Z => n7216);
   U5201 : IVI port map( A => n247, Z => n7217);
   U5202 : IVI port map( A => n247, Z => n7218);
   U5203 : IVI port map( A => n247, Z => n7219);
   U5204 : IVI port map( A => n247, Z => n7220);
   U5205 : IVI port map( A => n247, Z => n7221);
   U5206 : IVI port map( A => n247, Z => n7222);
   U5207 : IVI port map( A => n247, Z => n7223);
   U5208 : IVI port map( A => n247, Z => n7224);
   U5209 : IVI port map( A => n247, Z => n7225);
   U5210 : IVI port map( A => n247, Z => n7226);
   U5211 : IVI port map( A => n247, Z => n7227);
   U5212 : IVI port map( A => n247, Z => n7228);
   U5213 : IVI port map( A => n247, Z => n7229);
   U5214 : IVI port map( A => n247, Z => n7230);
   U5215 : IVI port map( A => n247, Z => n7231);
   U5216 : IVI port map( A => n247, Z => n7232);
   U5217 : IVI port map( A => n247, Z => n7233);
   U5218 : IVI port map( A => n7233, Z => n7236);
   U5219 : IVI port map( A => n244, Z => n7237);
   U5220 : IVI port map( A => n244, Z => n7238);
   U5221 : IVI port map( A => n244, Z => n7239);
   U5222 : IVI port map( A => n244, Z => n7240);
   U5223 : IVI port map( A => n244, Z => n7241);
   U5224 : IVI port map( A => n244, Z => n7242);
   U5225 : IVI port map( A => n244, Z => n7243);
   U5226 : IVI port map( A => n244, Z => n7244);
   U5227 : IVI port map( A => n244, Z => n7245);
   U5228 : IVI port map( A => n244, Z => n7246);
   U5229 : IVI port map( A => n244, Z => n7247);
   U5230 : IVI port map( A => n244, Z => n7248);
   U5231 : IVI port map( A => n244, Z => n7249);
   U5232 : IVI port map( A => n244, Z => n7250);
   U5233 : IVI port map( A => n244, Z => n7251);
   U5234 : IVI port map( A => n244, Z => n7252);
   U5235 : IVI port map( A => n244, Z => n7253);
   U5236 : IVI port map( A => n7253, Z => n7256);
   U5237 : IVI port map( A => n182, Z => n7257);
   U5238 : IVI port map( A => n182, Z => n7258);
   U5239 : IVI port map( A => n182, Z => n7259);
   U5240 : IVI port map( A => n182, Z => n7260);
   U5241 : IVI port map( A => n182, Z => n7261);
   U5242 : IVI port map( A => n182, Z => n7262);
   U5243 : IVI port map( A => n182, Z => n7263);
   U5244 : IVI port map( A => n182, Z => n7264);
   U5245 : IVI port map( A => n182, Z => n7265);
   U5246 : IVI port map( A => n182, Z => n7266);
   U5247 : IVI port map( A => n182, Z => n7267);
   U5248 : IVI port map( A => n182, Z => n7268);
   U5249 : IVI port map( A => n182, Z => n7269);
   U5250 : IVI port map( A => n182, Z => n7270);
   U5251 : IVI port map( A => n182, Z => n7271);
   U5252 : IVI port map( A => n182, Z => n7272);
   U5253 : IVI port map( A => n182, Z => n7273);
   U5254 : IVI port map( A => n7273, Z => n7276);
   U5255 : IVI port map( A => n181, Z => n7277);
   U5256 : IVI port map( A => n181, Z => n7278);
   U5257 : IVI port map( A => n181, Z => n7279);
   U5258 : IVI port map( A => n181, Z => n7280);
   U5259 : IVI port map( A => n181, Z => n7281);
   U5260 : IVI port map( A => n181, Z => n7282);
   U5261 : IVI port map( A => n181, Z => n7283);
   U5262 : IVI port map( A => n181, Z => n7284);
   U5263 : IVI port map( A => n181, Z => n7285);
   U5264 : IVI port map( A => n181, Z => n7286);
   U5265 : IVI port map( A => n181, Z => n7287);
   U5266 : IVI port map( A => n181, Z => n7288);
   U5267 : IVI port map( A => n181, Z => n7289);
   U5268 : IVI port map( A => n181, Z => n7290);
   U5269 : IVI port map( A => n181, Z => n7291);
   U5270 : IVI port map( A => n181, Z => n7292);
   U5271 : IVI port map( A => n181, Z => n7293);
   U5272 : IVI port map( A => n7293, Z => n7296);
   U5273 : IVI port map( A => n171, Z => n7297);
   U5274 : IVI port map( A => n171, Z => n7298);
   U5275 : IVI port map( A => n171, Z => n7299);
   U5276 : IVI port map( A => n171, Z => n7300);
   U5277 : IVI port map( A => n171, Z => n7301);
   U5278 : IVI port map( A => n171, Z => n7302);
   U5279 : IVI port map( A => n171, Z => n7303);
   U5280 : IVI port map( A => n171, Z => n7304);
   U5281 : IVI port map( A => n171, Z => n7305);
   U5282 : IVI port map( A => n171, Z => n7306);
   U5283 : IVI port map( A => n171, Z => n7307);
   U5284 : IVI port map( A => n171, Z => n7308);
   U5285 : IVI port map( A => n171, Z => n7309);
   U5286 : IVI port map( A => n171, Z => n7310);
   U5287 : IVI port map( A => n171, Z => n7311);
   U5288 : IVI port map( A => n171, Z => n7312);
   U5289 : IVI port map( A => n171, Z => n7313);
   U5290 : IVI port map( A => n7313, Z => n7316);
   U5291 : IVI port map( A => n170, Z => n7317);
   U5292 : IVI port map( A => n170, Z => n7318);
   U5293 : IVI port map( A => n170, Z => n7319);
   U5294 : IVI port map( A => n170, Z => n7320);
   U5295 : IVI port map( A => n170, Z => n7321);
   U5296 : IVI port map( A => n170, Z => n7322);
   U5297 : IVI port map( A => n170, Z => n7323);
   U5298 : IVI port map( A => n170, Z => n7324);
   U5299 : IVI port map( A => n170, Z => n7325);
   U5300 : IVI port map( A => n170, Z => n7326);
   U5301 : IVI port map( A => n170, Z => n7327);
   U5302 : IVI port map( A => n170, Z => n7328);
   U5303 : IVI port map( A => n170, Z => n7329);
   U5304 : IVI port map( A => n170, Z => n7330);
   U5305 : IVI port map( A => n170, Z => n7331);
   U5306 : IVI port map( A => n170, Z => n7332);
   U5307 : IVI port map( A => n170, Z => n7333);
   U5308 : IVI port map( A => n7333, Z => n7336);
   U5309 : IVI port map( A => n243, Z => n7337);
   U5310 : IVI port map( A => n243, Z => n7338);
   U5311 : IVI port map( A => n243, Z => n7339);
   U5312 : IVI port map( A => n243, Z => n7340);
   U5313 : IVI port map( A => n243, Z => n7341);
   U5314 : IVI port map( A => n243, Z => n7342);
   U5315 : IVI port map( A => n243, Z => n7343);
   U5316 : IVI port map( A => n243, Z => n7344);
   U5317 : IVI port map( A => n243, Z => n7345);
   U5318 : IVI port map( A => n243, Z => n7346);
   U5319 : IVI port map( A => n243, Z => n7347);
   U5320 : IVI port map( A => n243, Z => n7348);
   U5321 : IVI port map( A => n243, Z => n7349);
   U5322 : IVI port map( A => n243, Z => n7350);
   U5323 : IVI port map( A => n243, Z => n7351);
   U5324 : IVI port map( A => n243, Z => n7352);
   U5325 : IVI port map( A => n243, Z => n7353);
   U5326 : IVI port map( A => n7353, Z => n7356);
   U5327 : IVI port map( A => n242, Z => n7357);
   U5328 : IVI port map( A => n242, Z => n7358);
   U5329 : IVI port map( A => n242, Z => n7359);
   U5330 : IVI port map( A => n242, Z => n7360);
   U5331 : IVI port map( A => n242, Z => n7361);
   U5332 : IVI port map( A => n242, Z => n7362);
   U5333 : IVI port map( A => n242, Z => n7363);
   U5334 : IVI port map( A => n242, Z => n7364);
   U5335 : IVI port map( A => n242, Z => n7365);
   U5336 : IVI port map( A => n242, Z => n7366);
   U5337 : IVI port map( A => n242, Z => n7367);
   U5338 : IVI port map( A => n242, Z => n7368);
   U5339 : IVI port map( A => n242, Z => n7369);
   U5340 : IVI port map( A => n242, Z => n7370);
   U5341 : IVI port map( A => n242, Z => n7371);
   U5342 : IVI port map( A => n242, Z => n7372);
   U5343 : IVI port map( A => n242, Z => n7373);
   U5344 : IVI port map( A => n7373, Z => n7376);
   U5345 : IVI port map( A => n241, Z => n7377);
   U5346 : IVI port map( A => n241, Z => n7378);
   U5347 : IVI port map( A => n241, Z => n7379);
   U5348 : IVI port map( A => n241, Z => n7380);
   U5349 : IVI port map( A => n241, Z => n7381);
   U5350 : IVI port map( A => n241, Z => n7382);
   U5351 : IVI port map( A => n241, Z => n7383);
   U5352 : IVI port map( A => n241, Z => n7384);
   U5353 : IVI port map( A => n241, Z => n7385);
   U5354 : IVI port map( A => n241, Z => n7386);
   U5355 : IVI port map( A => n241, Z => n7387);
   U5356 : IVI port map( A => n241, Z => n7388);
   U5357 : IVI port map( A => n241, Z => n7389);
   U5358 : IVI port map( A => n241, Z => n7390);
   U5359 : IVI port map( A => n241, Z => n7391);
   U5360 : IVI port map( A => n241, Z => n7392);
   U5361 : IVI port map( A => n241, Z => n7393);
   U5362 : IVI port map( A => n7393, Z => n7396);
   U5363 : IVI port map( A => n240, Z => n7397);
   U5364 : IVI port map( A => n240, Z => n7398);
   U5365 : IVI port map( A => n240, Z => n7399);
   U5366 : IVI port map( A => n240, Z => n7400);
   U5367 : IVI port map( A => n240, Z => n7401);
   U5368 : IVI port map( A => n240, Z => n7402);
   U5369 : IVI port map( A => n240, Z => n7403);
   U5370 : IVI port map( A => n240, Z => n7404);
   U5371 : IVI port map( A => n240, Z => n7405);
   U5372 : IVI port map( A => n240, Z => n7406);
   U5373 : IVI port map( A => n240, Z => n7407);
   U5374 : IVI port map( A => n240, Z => n7408);
   U5375 : IVI port map( A => n240, Z => n7409);
   U5376 : IVI port map( A => n240, Z => n7410);
   U5377 : IVI port map( A => n240, Z => n7411);
   U5378 : IVI port map( A => n240, Z => n7412);
   U5379 : IVI port map( A => n240, Z => n7413);
   U5380 : IVI port map( A => n7413, Z => n7416);
   U5381 : IVI port map( A => n169, Z => n7417);
   U5382 : IVI port map( A => n169, Z => n7418);
   U5383 : IVI port map( A => n169, Z => n7419);
   U5384 : IVI port map( A => n169, Z => n7420);
   U5385 : IVI port map( A => n169, Z => n7421);
   U5386 : IVI port map( A => n169, Z => n7422);
   U5387 : IVI port map( A => n169, Z => n7423);
   U5388 : IVI port map( A => n169, Z => n7424);
   U5389 : IVI port map( A => n169, Z => n7425);
   U5390 : IVI port map( A => n169, Z => n7426);
   U5391 : IVI port map( A => n169, Z => n7427);
   U5392 : IVI port map( A => n169, Z => n7428);
   U5393 : IVI port map( A => n169, Z => n7429);
   U5394 : IVI port map( A => n169, Z => n7430);
   U5395 : IVI port map( A => n169, Z => n7431);
   U5396 : IVI port map( A => n169, Z => n7432);
   U5397 : IVI port map( A => n169, Z => n7433);
   U5398 : IVI port map( A => n7433, Z => n7436);
   U5399 : IVI port map( A => n163, Z => n7437);
   U5400 : IVI port map( A => n163, Z => n7438);
   U5401 : IVI port map( A => n163, Z => n7439);
   U5402 : IVI port map( A => n163, Z => n7440);
   U5403 : IVI port map( A => n163, Z => n7441);
   U5404 : IVI port map( A => n163, Z => n7442);
   U5405 : IVI port map( A => n163, Z => n7443);
   U5406 : IVI port map( A => n163, Z => n7444);
   U5407 : IVI port map( A => n163, Z => n7445);
   U5408 : IVI port map( A => n163, Z => n7446);
   U5409 : IVI port map( A => n163, Z => n7447);
   U5410 : IVI port map( A => n163, Z => n7448);
   U5411 : IVI port map( A => n163, Z => n7449);
   U5412 : IVI port map( A => n163, Z => n7450);
   U5413 : IVI port map( A => n163, Z => n7451);
   U5414 : IVI port map( A => n163, Z => n7452);
   U5415 : IVI port map( A => n163, Z => n7453);
   U5416 : IVI port map( A => n7453, Z => n7456);
   U5417 : IVI port map( A => n150, Z => n7457);
   U5418 : IVI port map( A => n150, Z => n7458);
   U5419 : IVI port map( A => n150, Z => n7459);
   U5420 : IVI port map( A => n150, Z => n7460);
   U5421 : IVI port map( A => n150, Z => n7461);
   U5422 : IVI port map( A => n150, Z => n7462);
   U5423 : IVI port map( A => n150, Z => n7463);
   U5424 : IVI port map( A => n150, Z => n7464);
   U5425 : IVI port map( A => n150, Z => n7465);
   U5426 : IVI port map( A => n150, Z => n7466);
   U5427 : IVI port map( A => n150, Z => n7467);
   U5428 : IVI port map( A => n150, Z => n7468);
   U5429 : IVI port map( A => n150, Z => n7469);
   U5430 : IVI port map( A => n150, Z => n7470);
   U5431 : IVI port map( A => n150, Z => n7471);
   U5432 : IVI port map( A => n150, Z => n7472);
   U5433 : IVI port map( A => n150, Z => n7473);
   U5434 : IVI port map( A => n7473, Z => n7476);
   U5435 : IVI port map( A => n122, Z => n7477);
   U5436 : IVI port map( A => n122, Z => n7478);
   U5437 : IVI port map( A => n122, Z => n7479);
   U5438 : IVI port map( A => n122, Z => n7480);
   U5439 : IVI port map( A => n122, Z => n7481);
   U5440 : IVI port map( A => n122, Z => n7482);
   U5441 : IVI port map( A => n122, Z => n7483);
   U5442 : IVI port map( A => n122, Z => n7484);
   U5443 : IVI port map( A => n122, Z => n7485);
   U5444 : IVI port map( A => n122, Z => n7486);
   U5445 : IVI port map( A => n122, Z => n7487);
   U5446 : IVI port map( A => n122, Z => n7488);
   U5447 : IVI port map( A => n122, Z => n7489);
   U5448 : IVI port map( A => n122, Z => n7490);
   U5449 : IVI port map( A => n122, Z => n7491);
   U5450 : IVI port map( A => n122, Z => n7492);
   U5451 : IVI port map( A => n122, Z => n7493);
   U5452 : IVI port map( A => n7493, Z => n7496);
   U5453 : IVI port map( A => n109, Z => n7497);
   U5454 : IVI port map( A => n109, Z => n7498);
   U5455 : IVI port map( A => n109, Z => n7499);
   U5456 : IVI port map( A => n109, Z => n7500);
   U5457 : IVI port map( A => n109, Z => n7501);
   U5458 : IVI port map( A => n109, Z => n7502);
   U5459 : IVI port map( A => n109, Z => n7503);
   U5460 : IVI port map( A => n109, Z => n7504);
   U5461 : IVI port map( A => n109, Z => n7505);
   U5462 : IVI port map( A => n109, Z => n7506);
   U5463 : IVI port map( A => n109, Z => n7507);
   U5464 : IVI port map( A => n109, Z => n7508);
   U5465 : IVI port map( A => n109, Z => n7509);
   U5466 : IVI port map( A => n109, Z => n7510);
   U5467 : IVI port map( A => n109, Z => n7511);
   U5468 : IVI port map( A => n109, Z => n7512);
   U5469 : IVI port map( A => n109, Z => n7513);
   U5470 : IVI port map( A => n7513, Z => n7516);
   U5471 : IVI port map( A => n81, Z => n7517);
   U5472 : IVI port map( A => n81, Z => n7518);
   U5473 : IVI port map( A => n81, Z => n7519);
   U5474 : IVI port map( A => n81, Z => n7520);
   U5475 : IVI port map( A => n81, Z => n7521);
   U5476 : IVI port map( A => n81, Z => n7522);
   U5477 : IVI port map( A => n81, Z => n7523);
   U5478 : IVI port map( A => n81, Z => n7524);
   U5479 : IVI port map( A => n81, Z => n7525);
   U5480 : IVI port map( A => n81, Z => n7526);
   U5481 : IVI port map( A => n81, Z => n7527);
   U5482 : IVI port map( A => n81, Z => n7528);
   U5483 : IVI port map( A => n81, Z => n7529);
   U5484 : IVI port map( A => n81, Z => n7530);
   U5485 : IVI port map( A => n81, Z => n7531);
   U5486 : IVI port map( A => n81, Z => n7532);
   U5487 : IVI port map( A => n81, Z => n7533);
   U5488 : IVI port map( A => n7533, Z => n7536);
   U5489 : IVI port map( A => n72, Z => n7537);
   U5490 : IVI port map( A => n72, Z => n7538);
   U5491 : IVI port map( A => n72, Z => n7539);
   U5492 : IVI port map( A => n72, Z => n7540);
   U5493 : IVI port map( A => n72, Z => n7541);
   U5494 : IVI port map( A => n72, Z => n7542);
   U5495 : IVI port map( A => n72, Z => n7543);
   U5496 : IVI port map( A => n72, Z => n7544);
   U5497 : IVI port map( A => n72, Z => n7545);
   U5498 : IVI port map( A => n72, Z => n7546);
   U5499 : IVI port map( A => n72, Z => n7547);
   U5500 : IVI port map( A => n72, Z => n7548);
   U5501 : IVI port map( A => n72, Z => n7549);
   U5502 : IVI port map( A => n72, Z => n7550);
   U5503 : IVI port map( A => n72, Z => n7551);
   U5504 : IVI port map( A => n72, Z => n7552);
   U5505 : IVI port map( A => n72, Z => n7553);
   U5506 : IVI port map( A => n7553, Z => n7556);
   U5507 : IVI port map( A => n71, Z => n7557);
   U5508 : IVI port map( A => n71, Z => n7558);
   U5509 : IVI port map( A => n71, Z => n7559);
   U5510 : IVI port map( A => n71, Z => n7560);
   U5511 : IVI port map( A => n71, Z => n7561);
   U5512 : IVI port map( A => n71, Z => n7562);
   U5513 : IVI port map( A => n71, Z => n7563);
   U5514 : IVI port map( A => n71, Z => n7564);
   U5515 : IVI port map( A => n71, Z => n7565);
   U5516 : IVI port map( A => n71, Z => n7566);
   U5517 : IVI port map( A => n71, Z => n7567);
   U5518 : IVI port map( A => n71, Z => n7568);
   U5519 : IVI port map( A => n71, Z => n7569);
   U5520 : IVI port map( A => n71, Z => n7570);
   U5521 : IVI port map( A => n71, Z => n7571);
   U5522 : IVI port map( A => n71, Z => n7572);
   U5523 : IVI port map( A => n71, Z => n7573);
   U5524 : IVI port map( A => n7573, Z => n7576);
   U5525 : IVI port map( A => n69, Z => n7577);
   U5526 : IVI port map( A => n69, Z => n7578);
   U5527 : IVI port map( A => n69, Z => n7579);
   U5528 : IVI port map( A => n69, Z => n7580);
   U5529 : IVI port map( A => n69, Z => n7581);
   U5530 : IVI port map( A => n69, Z => n7582);
   U5531 : IVI port map( A => n69, Z => n7583);
   U5532 : IVI port map( A => n69, Z => n7584);
   U5533 : IVI port map( A => n69, Z => n7585);
   U5534 : IVI port map( A => n69, Z => n7586);
   U5535 : IVI port map( A => n69, Z => n7587);
   U5536 : IVI port map( A => n69, Z => n7588);
   U5537 : IVI port map( A => n69, Z => n7589);
   U5538 : IVI port map( A => n69, Z => n7590);
   U5539 : IVI port map( A => n69, Z => n7591);
   U5540 : IVI port map( A => n69, Z => n7592);
   U5541 : IVI port map( A => n69, Z => n7593);
   U5542 : IVI port map( A => n7593, Z => n7596);
   U5543 : IVI port map( A => n63, Z => n7597);
   U5544 : IVI port map( A => n63, Z => n7598);
   U5545 : IVI port map( A => n63, Z => n7599);
   U5546 : IVI port map( A => n63, Z => n7600);
   U5547 : IVI port map( A => n63, Z => n7601);
   U5548 : IVI port map( A => n63, Z => n7602);
   U5549 : IVI port map( A => n63, Z => n7603);
   U5550 : IVI port map( A => n63, Z => n7604);
   U5551 : IVI port map( A => n63, Z => n7605);
   U5552 : IVI port map( A => n63, Z => n7606);
   U5553 : IVI port map( A => n63, Z => n7607);
   U5554 : IVI port map( A => n63, Z => n7608);
   U5555 : IVI port map( A => n63, Z => n7609);
   U5556 : IVI port map( A => n63, Z => n7610);
   U5557 : IVI port map( A => n63, Z => n7611);
   U5558 : IVI port map( A => n63, Z => n7612);
   U5559 : IVI port map( A => n63, Z => n7613);
   U5560 : IVI port map( A => n7613, Z => n7616);
   U5561 : IVI port map( A => n59, Z => n7617);
   U5562 : IVI port map( A => n59, Z => n7618);
   U5563 : IVI port map( A => n59, Z => n7619);
   U5564 : IVI port map( A => n59, Z => n7620);
   U5565 : IVI port map( A => n59, Z => n7621);
   U5566 : IVI port map( A => n59, Z => n7622);
   U5567 : IVI port map( A => n59, Z => n7623);
   U5568 : IVI port map( A => n59, Z => n7624);
   U5569 : IVI port map( A => n59, Z => n7625);
   U5570 : IVI port map( A => n59, Z => n7626);
   U5571 : IVI port map( A => n59, Z => n7627);
   U5572 : IVI port map( A => n59, Z => n7628);
   U5573 : IVI port map( A => n59, Z => n7629);
   U5574 : IVI port map( A => n59, Z => n7630);
   U5575 : IVI port map( A => n59, Z => n7631);
   U5576 : IVI port map( A => n59, Z => n7632);
   U5577 : IVI port map( A => n59, Z => n7633);
   U5578 : IVI port map( A => n7633, Z => n7636);
   U5579 : IVI port map( A => n53, Z => n7637);
   U5580 : IVI port map( A => n53, Z => n7638);
   U5581 : IVI port map( A => n53, Z => n7639);
   U5582 : IVI port map( A => n53, Z => n7640);
   U5583 : IVI port map( A => n53, Z => n7641);
   U5584 : IVI port map( A => n53, Z => n7642);
   U5585 : IVI port map( A => n53, Z => n7643);
   U5586 : IVI port map( A => n53, Z => n7644);
   U5587 : IVI port map( A => n53, Z => n7645);
   U5588 : IVI port map( A => n53, Z => n7646);
   U5589 : IVI port map( A => n53, Z => n7647);
   U5590 : IVI port map( A => n53, Z => n7648);
   U5591 : IVI port map( A => n53, Z => n7649);
   U5592 : IVI port map( A => n53, Z => n7650);
   U5593 : IVI port map( A => n53, Z => n7651);
   U5594 : IVI port map( A => n53, Z => n7652);
   U5595 : IVI port map( A => n53, Z => n7653);
   U5596 : IVI port map( A => n7653, Z => n7656);
   U5597 : IVI port map( A => n48, Z => n7657);
   U5598 : IVI port map( A => n48, Z => n7658);
   U5599 : IVI port map( A => n48, Z => n7659);
   U5600 : IVI port map( A => n48, Z => n7660);
   U5601 : IVI port map( A => n48, Z => n7661);
   U5602 : IVI port map( A => n48, Z => n7662);
   U5603 : IVI port map( A => n48, Z => n7663);
   U5604 : IVI port map( A => n48, Z => n7664);
   U5605 : IVI port map( A => n48, Z => n7665);
   U5606 : IVI port map( A => n48, Z => n7666);
   U5607 : IVI port map( A => n48, Z => n7667);
   U5608 : IVI port map( A => n48, Z => n7668);
   U5609 : IVI port map( A => n48, Z => n7669);
   U5610 : IVI port map( A => n48, Z => n7670);
   U5611 : IVI port map( A => n48, Z => n7671);
   U5612 : IVI port map( A => n48, Z => n7672);
   U5613 : IVI port map( A => n48, Z => n7673);
   U5614 : IVI port map( A => n7673, Z => n7676);
   U5615 : IVI port map( A => n43, Z => n7677);
   U5616 : IVI port map( A => n43, Z => n7678);
   U5617 : IVI port map( A => n43, Z => n7679);
   U5618 : IVI port map( A => n43, Z => n7680);
   U5619 : IVI port map( A => n43, Z => n7681);
   U5620 : IVI port map( A => n43, Z => n7682);
   U5621 : IVI port map( A => n43, Z => n7683);
   U5622 : IVI port map( A => n43, Z => n7684);
   U5623 : IVI port map( A => n43, Z => n7685);
   U5624 : IVI port map( A => n43, Z => n7686);
   U5625 : IVI port map( A => n43, Z => n7687);
   U5626 : IVI port map( A => n43, Z => n7688);
   U5627 : IVI port map( A => n43, Z => n7689);
   U5628 : IVI port map( A => n43, Z => n7690);
   U5629 : IVI port map( A => n43, Z => n7691);
   U5630 : IVI port map( A => n43, Z => n7692);
   U5631 : IVI port map( A => n43, Z => n7693);
   U5632 : IVI port map( A => n7693, Z => n7696);
   U5633 : IVI port map( A => n38, Z => n7697);
   U5634 : IVI port map( A => n38, Z => n7698);
   U5635 : IVI port map( A => n38, Z => n7699);
   U5636 : IVI port map( A => n38, Z => n7700);
   U5637 : IVI port map( A => n38, Z => n7701);
   U5638 : IVI port map( A => n38, Z => n7702);
   U5639 : IVI port map( A => n38, Z => n7703);
   U5640 : IVI port map( A => n38, Z => n7704);
   U5641 : IVI port map( A => n38, Z => n7705);
   U5642 : IVI port map( A => n38, Z => n7706);
   U5643 : IVI port map( A => n38, Z => n7707);
   U5644 : IVI port map( A => n38, Z => n7708);
   U5645 : IVI port map( A => n38, Z => n7709);
   U5646 : IVI port map( A => n38, Z => n7710);
   U5647 : IVI port map( A => n38, Z => n7711);
   U5648 : IVI port map( A => n38, Z => n7712);
   U5649 : IVI port map( A => n38, Z => n7713);
   U5650 : IVI port map( A => n7713, Z => n7716);
   U5651 : IVI port map( A => n33, Z => n7717);
   U5652 : IVI port map( A => n33, Z => n7718);
   U5653 : IVI port map( A => n33, Z => n7719);
   U5654 : IVI port map( A => n33, Z => n7720);
   U5655 : IVI port map( A => n33, Z => n7721);
   U5656 : IVI port map( A => n33, Z => n7722);
   U5657 : IVI port map( A => n33, Z => n7723);
   U5658 : IVI port map( A => n33, Z => n7724);
   U5659 : IVI port map( A => n33, Z => n7725);
   U5660 : IVI port map( A => n33, Z => n7726);
   U5661 : IVI port map( A => n33, Z => n7727);
   U5662 : IVI port map( A => n33, Z => n7728);
   U5663 : IVI port map( A => n33, Z => n7729);
   U5664 : IVI port map( A => n33, Z => n7730);
   U5665 : IVI port map( A => n33, Z => n7731);
   U5666 : IVI port map( A => n33, Z => n7732);
   U5667 : IVI port map( A => n33, Z => n7733);
   U5668 : IVI port map( A => n7733, Z => n7736);
   U5669 : IVI port map( A => n28, Z => n7737);
   U5670 : IVI port map( A => n28, Z => n7738);
   U5671 : IVI port map( A => n28, Z => n7739);
   U5672 : IVI port map( A => n28, Z => n7740);
   U5673 : IVI port map( A => n28, Z => n7741);
   U5674 : IVI port map( A => n28, Z => n7742);
   U5675 : IVI port map( A => n28, Z => n7743);
   U5676 : IVI port map( A => n28, Z => n7744);
   U5677 : IVI port map( A => n28, Z => n7745);
   U5678 : IVI port map( A => n28, Z => n7746);
   U5679 : IVI port map( A => n28, Z => n7747);
   U5680 : IVI port map( A => n28, Z => n7748);
   U5681 : IVI port map( A => n28, Z => n7749);
   U5682 : IVI port map( A => n28, Z => n7750);
   U5683 : IVI port map( A => n28, Z => n7751);
   U5684 : IVI port map( A => n28, Z => n7752);
   U5685 : IVI port map( A => n28, Z => n7753);
   U5686 : IVI port map( A => n7753, Z => n7756);
   U5687 : IVI port map( A => n23, Z => n7757);
   U5688 : IVI port map( A => n23, Z => n7758);
   U5689 : IVI port map( A => n23, Z => n7759);
   U5690 : IVI port map( A => n23, Z => n7760);
   U5691 : IVI port map( A => n23, Z => n7761);
   U5692 : IVI port map( A => n23, Z => n7762);
   U5693 : IVI port map( A => n23, Z => n7763);
   U5694 : IVI port map( A => n23, Z => n7764);
   U5695 : IVI port map( A => n23, Z => n7765);
   U5696 : IVI port map( A => n23, Z => n7766);
   U5697 : IVI port map( A => n23, Z => n7767);
   U5698 : IVI port map( A => n23, Z => n7768);
   U5699 : IVI port map( A => n23, Z => n7769);
   U5700 : IVI port map( A => n23, Z => n7770);
   U5701 : IVI port map( A => n23, Z => n7771);
   U5702 : IVI port map( A => n23, Z => n7772);
   U5703 : IVI port map( A => n23, Z => n7773);
   U5704 : IVI port map( A => n7773, Z => n7776);
   U5705 : IVI port map( A => n22, Z => n7777);
   U5706 : IVI port map( A => n22, Z => n7778);
   U5707 : IVI port map( A => n22, Z => n7779);
   U5708 : IVI port map( A => n22, Z => n7780);
   U5709 : IVI port map( A => n22, Z => n7781);
   U5710 : IVI port map( A => n22, Z => n7782);
   U5711 : IVI port map( A => n22, Z => n7783);
   U5712 : IVI port map( A => n22, Z => n7784);
   U5713 : IVI port map( A => n22, Z => n7785);
   U5714 : IVI port map( A => n22, Z => n7786);
   U5715 : IVI port map( A => n22, Z => n7787);
   U5716 : IVI port map( A => n22, Z => n7788);
   U5717 : IVI port map( A => n22, Z => n7789);
   U5718 : IVI port map( A => n22, Z => n7790);
   U5719 : IVI port map( A => n22, Z => n7791);
   U5720 : IVI port map( A => n22, Z => n7792);
   U5721 : IVI port map( A => n22, Z => n7793);
   U5722 : IVI port map( A => n7793, Z => n7796);
   U5723 : IVI port map( A => n14, Z => n7797);
   U5724 : IVI port map( A => n14, Z => n7798);
   U5725 : IVI port map( A => n14, Z => n7799);
   U5726 : IVI port map( A => n14, Z => n7800);
   U5727 : IVI port map( A => n14, Z => n7801);
   U5728 : IVI port map( A => n14, Z => n7802);
   U5729 : IVI port map( A => n14, Z => n7803);
   U5730 : IVI port map( A => n14, Z => n7804);
   U5731 : IVI port map( A => n14, Z => n7805);
   U5732 : IVI port map( A => n14, Z => n7806);
   U5733 : IVI port map( A => n14, Z => n7807);
   U5734 : IVI port map( A => n14, Z => n7808);
   U5735 : IVI port map( A => n14, Z => n7809);
   U5736 : IVI port map( A => n14, Z => n7810);
   U5737 : IVI port map( A => n14, Z => n7811);
   U5738 : IVI port map( A => n14, Z => n7812);
   U5739 : IVI port map( A => n14, Z => n7813);
   U5740 : IVI port map( A => n7813, Z => n7816);
   U5741 : IVI port map( A => n12, Z => n7817);
   U5742 : IVI port map( A => n12, Z => n7818);
   U5743 : IVI port map( A => n12, Z => n7819);
   U5744 : IVI port map( A => n12, Z => n7820);
   U5745 : IVI port map( A => n12, Z => n7821);
   U5746 : IVI port map( A => n12, Z => n7822);
   U5747 : IVI port map( A => n12, Z => n7823);
   U5748 : IVI port map( A => n12, Z => n7824);
   U5749 : IVI port map( A => n12, Z => n7825);
   U5750 : IVI port map( A => n12, Z => n7826);
   U5751 : IVI port map( A => n12, Z => n7827);
   U5752 : IVI port map( A => n12, Z => n7828);
   U5753 : IVI port map( A => n12, Z => n7829);
   U5754 : IVI port map( A => n12, Z => n7830);
   U5755 : IVI port map( A => n12, Z => n7831);
   U5756 : IVI port map( A => n12, Z => n7832);
   U5757 : IVI port map( A => n12, Z => n7833);
   U5758 : IVI port map( A => n7833, Z => n7836);
   U5759 : IVI port map( A => n11, Z => n7837);
   U5760 : IVI port map( A => n11, Z => n7838);
   U5761 : IVI port map( A => n11, Z => n7839);
   U5762 : IVI port map( A => n11, Z => n7840);
   U5763 : IVI port map( A => n11, Z => n7841);
   U5764 : IVI port map( A => n11, Z => n7842);
   U5765 : IVI port map( A => n11, Z => n7843);
   U5766 : IVI port map( A => n11, Z => n7844);
   U5767 : IVI port map( A => n11, Z => n7845);
   U5768 : IVI port map( A => n11, Z => n7846);
   U5769 : IVI port map( A => n11, Z => n7847);
   U5770 : IVI port map( A => n11, Z => n7848);
   U5771 : IVI port map( A => n11, Z => n7849);
   U5772 : IVI port map( A => n11, Z => n7850);
   U5773 : IVI port map( A => n11, Z => n7851);
   U5774 : IVI port map( A => n11, Z => n7852);
   U5775 : IVI port map( A => n11, Z => n7853);
   U5776 : IVI port map( A => n7853, Z => n7856);
   U5777 : IVI port map( A => n10, Z => n7857);
   U5778 : IVI port map( A => n10, Z => n7858);
   U5779 : IVI port map( A => n10, Z => n7859);
   U5780 : IVI port map( A => n10, Z => n7860);
   U5781 : IVI port map( A => n10, Z => n7861);
   U5782 : IVI port map( A => n10, Z => n7862);
   U5783 : IVI port map( A => n10, Z => n7863);
   U5784 : IVI port map( A => n10, Z => n7864);
   U5785 : IVI port map( A => n10, Z => n7865);
   U5786 : IVI port map( A => n10, Z => n7866);
   U5787 : IVI port map( A => n10, Z => n7867);
   U5788 : IVI port map( A => n10, Z => n7868);
   U5789 : IVI port map( A => n10, Z => n7869);
   U5790 : IVI port map( A => n10, Z => n7870);
   U5791 : IVI port map( A => n10, Z => n7871);
   U5792 : IVI port map( A => n10, Z => n7872);
   U5793 : IVI port map( A => n10, Z => n7873);
   U5794 : IVI port map( A => n7873, Z => n7876);
   U5795 : IVI port map( A => n9, Z => n7877);
   U5796 : IVI port map( A => n9, Z => n7878);
   U5797 : IVI port map( A => n9, Z => n7879);
   U5798 : IVI port map( A => n9, Z => n7880);
   U5799 : IVI port map( A => n9, Z => n7881);
   U5800 : IVI port map( A => n9, Z => n7882);
   U5801 : IVI port map( A => n9, Z => n7883);
   U5802 : IVI port map( A => n9, Z => n7884);
   U5803 : IVI port map( A => n9, Z => n7885);
   U5804 : IVI port map( A => n9, Z => n7886);
   U5805 : IVI port map( A => n9, Z => n7887);
   U5806 : IVI port map( A => n9, Z => n7888);
   U5807 : IVI port map( A => n9, Z => n7889);
   U5808 : IVI port map( A => n9, Z => n7890);
   U5809 : IVI port map( A => n9, Z => n7891);
   U5810 : IVI port map( A => n9, Z => n7892);
   U5811 : IVI port map( A => n9, Z => n7893);
   U5812 : IVI port map( A => n7893, Z => n7896);
   U5813 : IVI port map( A => n8, Z => n7897);
   U5814 : IVI port map( A => n8, Z => n7898);
   U5815 : IVI port map( A => n8, Z => n7899);
   U5816 : IVI port map( A => n8, Z => n7900);
   U5817 : IVI port map( A => n8, Z => n7901);
   U5818 : IVI port map( A => n8, Z => n7902);
   U5819 : IVI port map( A => n8, Z => n7903);
   U5820 : IVI port map( A => n8, Z => n7904);
   U5821 : IVI port map( A => n8, Z => n7905);
   U5822 : IVI port map( A => n8, Z => n7906);
   U5823 : IVI port map( A => n8, Z => n7907);
   U5824 : IVI port map( A => n8, Z => n7908);
   U5825 : IVI port map( A => n8, Z => n7909);
   U5826 : IVI port map( A => n8, Z => n7910);
   U5827 : IVI port map( A => n8, Z => n7911);
   U5828 : IVI port map( A => n8, Z => n7912);
   U5829 : IVI port map( A => n8, Z => n7913);
   U5830 : IVI port map( A => n7913, Z => n7916);
   U5831 : IVI port map( A => n7, Z => n7917);
   U5832 : IVI port map( A => n7, Z => n7918);
   U5833 : IVI port map( A => n7, Z => n7919);
   U5834 : IVI port map( A => n7, Z => n7920);
   U5835 : IVI port map( A => n7, Z => n7921);
   U5836 : IVI port map( A => n7, Z => n7922);
   U5837 : IVI port map( A => n7, Z => n7923);
   U5838 : IVI port map( A => n7, Z => n7924);
   U5839 : IVI port map( A => n7, Z => n7925);
   U5840 : IVI port map( A => n7, Z => n7926);
   U5841 : IVI port map( A => n7, Z => n7927);
   U5842 : IVI port map( A => n7, Z => n7928);
   U5843 : IVI port map( A => n7, Z => n7929);
   U5844 : IVI port map( A => n7, Z => n7930);
   U5845 : IVI port map( A => n7, Z => n7931);
   U5846 : IVI port map( A => n7, Z => n7932);
   U5847 : IVI port map( A => n7, Z => n7933);
   U5848 : IVI port map( A => n7933, Z => n7936);
   U5849 : IVI port map( A => n6, Z => n7937);
   U5850 : IVI port map( A => n6, Z => n7938);
   U5851 : IVI port map( A => n6, Z => n7939);
   U5852 : IVI port map( A => n6, Z => n7940);
   U5853 : IVI port map( A => n6, Z => n7941);
   U5854 : IVI port map( A => n6, Z => n7942);
   U5855 : IVI port map( A => n6, Z => n7943);
   U5856 : IVI port map( A => n6, Z => n7944);
   U5857 : IVI port map( A => n6, Z => n7945);
   U5858 : IVI port map( A => n6, Z => n7946);
   U5859 : IVI port map( A => n6, Z => n7947);
   U5860 : IVI port map( A => n6, Z => n7948);
   U5861 : IVI port map( A => n6, Z => n7949);
   U5862 : IVI port map( A => n6, Z => n7950);
   U5863 : IVI port map( A => n6, Z => n7951);
   U5864 : IVI port map( A => n6, Z => n7952);
   U5865 : IVI port map( A => n6, Z => n7953);
   U5866 : IVI port map( A => n7953, Z => n7956);
   U5867 : IVI port map( A => n5, Z => n7957);
   U5868 : IVI port map( A => n5, Z => n7958);
   U5869 : IVI port map( A => n5, Z => n7959);
   U5870 : IVI port map( A => n5, Z => n7960);
   U5871 : IVI port map( A => n5, Z => n7961);
   U5872 : IVI port map( A => n5, Z => n7962);
   U5873 : IVI port map( A => n5, Z => n7963);
   U5874 : IVI port map( A => n5, Z => n7964);
   U5875 : IVI port map( A => n5, Z => n7965);
   U5876 : IVI port map( A => n5, Z => n7966);
   U5877 : IVI port map( A => n5, Z => n7967);
   U5878 : IVI port map( A => n5, Z => n7968);
   U5879 : IVI port map( A => n5, Z => n7969);
   U5880 : IVI port map( A => n5, Z => n7970);
   U5881 : IVI port map( A => n5, Z => n7971);
   U5882 : IVI port map( A => n5, Z => n7972);
   U5883 : IVI port map( A => n5, Z => n7973);
   U5884 : IVI port map( A => n7973, Z => n7976);
   U5885 : IVI port map( A => n4, Z => n7977);
   U5886 : IVI port map( A => n4, Z => n7978);
   U5887 : IVI port map( A => n4, Z => n7979);
   U5888 : IVI port map( A => n4, Z => n7980);
   U5889 : IVI port map( A => n4, Z => n7981);
   U5890 : IVI port map( A => n4, Z => n7982);
   U5891 : IVI port map( A => n4, Z => n7983);
   U5892 : IVI port map( A => n4, Z => n7984);
   U5893 : IVI port map( A => n4, Z => n7985);
   U5894 : IVI port map( A => n4, Z => n7986);
   U5895 : IVI port map( A => n4, Z => n7987);
   U5896 : IVI port map( A => n4, Z => n7988);
   U5897 : IVI port map( A => n4, Z => n7989);
   U5898 : IVI port map( A => n4, Z => n7990);
   U5899 : IVI port map( A => n4, Z => n7991);
   U5900 : IVI port map( A => n4, Z => n7992);
   U5901 : IVI port map( A => n4, Z => n7993);
   U5902 : IVI port map( A => n7993, Z => n7996);
   U5903 : IVI port map( A => n3, Z => n7997);
   U5904 : IVI port map( A => n3, Z => n7998);
   U5905 : IVI port map( A => n3, Z => n7999);
   U5906 : IVI port map( A => n3, Z => n8000);
   U5907 : IVI port map( A => n3, Z => n8001);
   U5908 : IVI port map( A => n3, Z => n8002);
   U5909 : IVI port map( A => n3, Z => n8003);
   U5910 : IVI port map( A => n3, Z => n8004);
   U5911 : IVI port map( A => n3, Z => n8005);
   U5912 : IVI port map( A => n3, Z => n8006);
   U5913 : IVI port map( A => n3, Z => n8007);
   U5914 : IVI port map( A => n3, Z => n8008);
   U5915 : IVI port map( A => n3, Z => n8009);
   U5916 : IVI port map( A => n3, Z => n8010);
   U5917 : IVI port map( A => n3, Z => n8011);
   U5918 : IVI port map( A => n3, Z => n8012);
   U5919 : IVI port map( A => n3, Z => n8013);
   U5920 : IVI port map( A => n8013, Z => n8016);
   U5921 : IVI port map( A => n2, Z => n8017);
   U5922 : IVI port map( A => n2, Z => n8018);
   U5923 : IVI port map( A => n2, Z => n8019);
   U5924 : IVI port map( A => n2, Z => n8020);
   U5925 : IVI port map( A => n2, Z => n8021);
   U5926 : IVI port map( A => n2, Z => n8022);
   U5927 : IVI port map( A => n2, Z => n8023);
   U5928 : IVI port map( A => n2, Z => n8024);
   U5929 : IVI port map( A => n2, Z => n8025);
   U5930 : IVI port map( A => n2, Z => n8026);
   U5931 : IVI port map( A => n2, Z => n8027);
   U5932 : IVI port map( A => n2, Z => n8028);
   U5933 : IVI port map( A => n2, Z => n8029);
   U5934 : IVI port map( A => n2, Z => n8030);
   U5935 : IVI port map( A => n2, Z => n8031);
   U5936 : IVI port map( A => n2, Z => n8032);
   U5937 : IVI port map( A => n2, Z => n8033);
   U5938 : IVI port map( A => n8033, Z => n8036);
   U5939 : IVI port map( A => n1, Z => n8037);
   U5940 : IVI port map( A => n1, Z => n8038);
   U5941 : IVI port map( A => n1, Z => n8039);
   U5942 : IVI port map( A => n1, Z => n8040);
   U5943 : IVI port map( A => n1, Z => n8041);
   U5944 : IVI port map( A => n1, Z => n8042);
   U5945 : IVI port map( A => n1, Z => n8043);
   U5946 : IVI port map( A => n1, Z => n8044);
   U5947 : IVI port map( A => n1, Z => n8045);
   U5948 : IVI port map( A => n1, Z => n8046);
   U5949 : IVI port map( A => n1, Z => n8047);
   U5950 : IVI port map( A => n1, Z => n8048);
   U5951 : IVI port map( A => n1, Z => n8049);
   U5952 : IVI port map( A => n1, Z => n8050);
   U5953 : IVI port map( A => n1, Z => n8051);
   U5954 : IVI port map( A => n1, Z => n8052);
   U5955 : IVI port map( A => n1, Z => n8053);
   U5956 : IVI port map( A => n8053, Z => n8056);
   U5957 : IVI port map( A => n8062, Z => n8061);
   U5958 : IVI port map( A => n2291, Z => n8062);
   U5959 : IVI port map( A => n444, Z => n8063);
   U5960 : IVI port map( A => n1883, Z => n8064);
   U5961 : IVI port map( A => n445, Z => n8065);
   U5962 : IVI port map( A => n446, Z => n8066);
   U5963 : IVI port map( A => n447, Z => n8067);
   U5964 : IVI port map( A => n1885, Z => n8068);
   U5965 : IVI port map( A => n1279, Z => n8069);
   U5966 : IVI port map( A => n1323, Z => n8070);
   U5967 : IVI port map( A => n440, Z => n8071);
   U5968 : IVI port map( A => n1864, Z => n8072);
   U5969 : IVI port map( A => n441, Z => n8073);
   U5970 : IVI port map( A => n442, Z => n8074);
   U5971 : IVI port map( A => n443, Z => n8075);
   U5972 : IVI port map( A => n1865, Z => n8076);
   U5973 : IVI port map( A => n1148, Z => n8077);
   U5974 : IVI port map( A => n1192, Z => n8078);
   U5975 : IVI port map( A => n432, Z => n8079);
   U5976 : IVI port map( A => n1852, Z => n8080);
   U5977 : IVI port map( A => n433, Z => n8081);
   U5978 : IVI port map( A => n434, Z => n8082);
   U5979 : IVI port map( A => n439, Z => n8083);
   U5980 : IVI port map( A => n1862, Z => n8084);
   U5981 : IVI port map( A => n1017, Z => n8085);
   U5982 : IVI port map( A => n1104, Z => n8086);
   U5983 : IVI port map( A => n428, Z => n8087);
   U5984 : IVI port map( A => n1845, Z => n8088);
   U5985 : IVI port map( A => n429, Z => n8089);
   U5986 : IVI port map( A => n430, Z => n8090);
   U5987 : IVI port map( A => n431, Z => n8091);
   U5988 : IVI port map( A => n1848, Z => n8092);
   U5989 : IVI port map( A => n929, Z => n8093);
   U5990 : IVI port map( A => n973, Z => n8094);
   U5991 : IVI port map( A => n420, Z => n8095);
   U5992 : IVI port map( A => n1841, Z => n8096);
   U5993 : IVI port map( A => n421, Z => n8097);
   U5994 : IVI port map( A => n422, Z => n8098);
   U5995 : IVI port map( A => n427, Z => n8099);
   U5996 : IVI port map( A => n1842, Z => n8100);
   U5997 : IVI port map( A => n798, Z => n8101);
   U5998 : IVI port map( A => n842, Z => n8102);
   U5999 : IVI port map( A => n416, Z => n8103);
   U6000 : IVI port map( A => n1830, Z => n8104);
   U6001 : IVI port map( A => n417, Z => n8105);
   U6002 : IVI port map( A => n418, Z => n8106);
   U6003 : IVI port map( A => n419, Z => n8107);
   U6004 : IVI port map( A => n1831, Z => n8108);
   U6005 : IVI port map( A => n667, Z => n8109);
   U6006 : IVI port map( A => n754, Z => n8110);
   U6007 : IVI port map( A => n408, Z => n8111);
   U6008 : IVI port map( A => n1790, Z => n8112);
   U6009 : IVI port map( A => n409, Z => n8113);
   U6010 : IVI port map( A => n410, Z => n8114);
   U6011 : IVI port map( A => n415, Z => n8115);
   U6012 : IVI port map( A => n1791, Z => n8116);
   U6013 : IVI port map( A => n579, Z => n8117);
   U6014 : IVI port map( A => n623, Z => n8118);
   U6015 : IVI port map( A => n404, Z => n8119);
   U6016 : IVI port map( A => n1674, Z => n8120);
   U6017 : IVI port map( A => n405, Z => n8121);
   U6018 : IVI port map( A => n406, Z => n8122);
   U6019 : IVI port map( A => n407, Z => n8123);
   U6020 : IVI port map( A => n1718, Z => n8124);
   U6021 : IVI port map( A => n491, Z => n8125);
   U6022 : IVI port map( A => n535, Z => n8126);
   U6023 : IVI port map( A => n8137, Z => n8127);
   U6024 : IVI port map( A => n8137, Z => n8128);
   U6025 : IVI port map( A => n8136, Z => n8129);
   U6026 : IVI port map( A => n8136, Z => n8130);
   U6027 : IVI port map( A => n8136, Z => n8131);
   U6028 : IVI port map( A => n8135, Z => n8132);
   U6029 : IVI port map( A => n8135, Z => n8133);
   U6030 : IVI port map( A => n8135, Z => n8134);
   U6031 : IVI port map( A => n8138, Z => n8135);
   U6032 : IVI port map( A => n8138, Z => n8136);
   U6033 : IVI port map( A => n8138, Z => n8137);
   U6034 : IVI port map( A => n8139, Z => n8138);
   U6035 : IVI port map( A => CE_I, Z => n8139);
   U6036 : IVI port map( A => n8166, Z => n8143);
   U6037 : IVI port map( A => n8127, Z => n8144);
   U6038 : IVI port map( A => n8127, Z => n8145);
   U6039 : IVI port map( A => n8127, Z => n8146);
   U6040 : IVI port map( A => n8128, Z => n8147);
   U6041 : IVI port map( A => n8128, Z => n8148);
   U6042 : IVI port map( A => n8128, Z => n8149);
   U6043 : IVI port map( A => n8129, Z => n8150);
   U6044 : IVI port map( A => n8129, Z => n8151);
   U6045 : IVI port map( A => n8129, Z => n8152);
   U6046 : IVI port map( A => n8130, Z => n8153);
   U6047 : IVI port map( A => n8130, Z => n8154);
   U6048 : IVI port map( A => n8130, Z => n8155);
   U6049 : IVI port map( A => n8131, Z => n8156);
   U6050 : IVI port map( A => n8131, Z => n8157);
   U6051 : IVI port map( A => n8131, Z => n8158);
   U6052 : IVI port map( A => n8132, Z => n8159);
   U6053 : IVI port map( A => n8132, Z => n8160);
   U6054 : IVI port map( A => n8132, Z => n8161);
   U6055 : IVI port map( A => n8133, Z => n8162);
   U6056 : IVI port map( A => n8133, Z => n8163);
   U6057 : IVI port map( A => n8133, Z => n8164);
   U6058 : IVI port map( A => n8134, Z => n8165);
   U6059 : IVI port map( A => n8134, Z => n8166);
   U6060 : ND2 port map( A => i_INTERN_ADDR_RD0_1_port, B => 
                           i_INTERN_ADDR_RD0_0_port, Z => n8167);
   U6061 : AN3 port map( A => i_INTERN_ADDR_RD0_1_port, B => 
                           i_INTERN_ADDR_RD0_0_port, C => 
                           i_INTERN_ADDR_RD0_2_port, Z => n8168);
   U6062 : ND2 port map( A => i_INTERN_ADDR_RD0_3_port, B => n8168, Z => n8169)
                           ;
   U6063 : NR2 port map( A => n8169, B => n6645, Z => n8170);
   U6064 : ND2 port map( A => i_SRAM_ADDR_WR0_1_port, B => 
                           i_SRAM_ADDR_WR0_0_port, Z => n8171);
   U6065 : AN3 port map( A => i_SRAM_ADDR_WR0_1_port, B => 
                           i_SRAM_ADDR_WR0_0_port, C => i_SRAM_ADDR_WR0_2_port,
                           Z => n8172);
   U6066 : ND2 port map( A => i_SRAM_ADDR_WR0_3_port, B => n8172, Z => n8173);
   U6067 : NR2 port map( A => n8173, B => n6639, Z => n8174);
   U6068 : ND2 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n8175);
   U6069 : EN port map( A => n8175, B => n2305, Z => N1749);
   U6070 : AN3 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, C => n2305, Z => n8177);
   U6071 : EO port map( A => n8177, B => v_CALCULATION_CNTR_3_port, Z => N1750)
                           ;
   U6072 : ND2 port map( A => v_CALCULATION_CNTR_3_port, B => n8177, Z => n8176
                           );
   U6073 : EN port map( A => n8176, B => v_CALCULATION_CNTR_4_port, Z => N1751)
                           ;
   U6074 : AN3 port map( A => v_CALCULATION_CNTR_3_port, B => n8177, C => 
                           v_CALCULATION_CNTR_4_port, Z => n8178);
   U6075 : EO port map( A => n8178, B => v_CALCULATION_CNTR_5_port, Z => N1752)
                           ;
   U6076 : ND2 port map( A => v_CALCULATION_CNTR_5_port, B => n8178, Z => n8179
                           );
   U6077 : EN port map( A => n8179, B => v_CALCULATION_CNTR_6_port, Z => N1753)
                           ;
   U6078 : NR2 port map( A => n8179, B => n2125, Z => n8180);
   U6079 : EO port map( A => v_CALCULATION_CNTR_7_port, B => n8180, Z => N1754)
                           ;
   U6080 : IVI port map( A => n326, Z => n8181);
   U6081 : IVI port map( A => n329, Z => n8182);
   U6082 : IVI port map( A => n330, Z => n8183);
   U6083 : IVI port map( A => n331, Z => n8184);
   U6084 : IVI port map( A => n332, Z => n8185);
   U6085 : IVI port map( A => n333, Z => n8186);
   U6086 : IVI port map( A => n334, Z => n8187);
   U6087 : IVI port map( A => n335, Z => n8188);
   U6088 : IVI port map( A => n328, Z => n8189);
   U6089 : IVI port map( A => n295, Z => n8190);
   U6090 : IVI port map( A => n298, Z => n8191);
   U6091 : IVI port map( A => n299, Z => n8192);
   U6092 : IVI port map( A => n300, Z => n8193);
   U6093 : IVI port map( A => n301, Z => n8194);
   U6094 : IVI port map( A => n302, Z => n8195);
   U6095 : IVI port map( A => n303, Z => n8196);
   U6096 : IVI port map( A => n304, Z => n8197);
   U6097 : IVI port map( A => n316, Z => n8198);
   U6098 : IVI port map( A => n319, Z => n8199);
   U6099 : IVI port map( A => n320, Z => n8200);
   U6100 : IVI port map( A => n321, Z => n8201);
   U6101 : IVI port map( A => n322, Z => n8202);
   U6102 : IVI port map( A => n323, Z => n8203);
   U6103 : IVI port map( A => n324, Z => n8204);
   U6104 : IVI port map( A => n325, Z => n8205);
   U6105 : IVI port map( A => n318, Z => n8206);
   U6106 : IVI port map( A => n305, Z => n8207);
   U6107 : IVI port map( A => n308, Z => n8208);
   U6108 : IVI port map( A => n309, Z => n8209);
   U6109 : IVI port map( A => n310, Z => n8210);
   U6110 : IVI port map( A => n311, Z => n8211);
   U6111 : IVI port map( A => n312, Z => n8212);
   U6112 : IVI port map( A => n313, Z => n8213);
   U6113 : IVI port map( A => n314, Z => n8214);
   U6114 : IVI port map( A => n283, Z => n8215);
   U6115 : IVI port map( A => n272, Z => n8216);
   U6116 : IVI port map( A => n2484, Z => n8217);
   U6117 : IVI port map( A => n2485, Z => n8218);
   U6118 : IVI port map( A => n2486, Z => n8219);
   U6119 : IVI port map( A => n57, Z => n8220);
   U6120 : IVI port map( A => n64, Z => n8221);
   U6121 : IVI port map( A => n2044, Z => n8222);
   U6122 : IVI port map( A => n1995, Z => n8223);
   U6123 : IVI port map( A => n1882, Z => n8224);
   U6124 : IVI port map( A => n2263, Z => n8225);
   U6125 : IVI port map( A => n2127, Z => n8226);
   U6126 : IVI port map( A => n1922, Z => n8227);
   U6127 : IVI port map( A => n2010, Z => n8228);
   U6128 : IVI port map( A => n1973, Z => n8229);
   U6129 : IVI port map( A => n2082, Z => n8230);
   U6130 : IVI port map( A => n1857, Z => n8231);
   U6131 : IVI port map( A => n2088, Z => n8232);
   U6132 : IVI port map( A => n2147, Z => n8233);
   U6133 : IVI port map( A => n2167, Z => n8234);
   U6134 : IVI port map( A => n2104, Z => n8235);
   U6135 : IVI port map( A => n1872, Z => n8237);
   U6136 : IVI port map( A => n2089, Z => n8238);
   U6137 : IVI port map( A => n1994, Z => n8239);
   U6138 : IVI port map( A => n2128, Z => n8240);
   U6139 : IVI port map( A => n1928, Z => n8241);
   U6140 : IVI port map( A => n2054, Z => n8242);
   U6141 : IVI port map( A => n2065, Z => n8243);
   U6142 : IVI port map( A => n2011, Z => n8244);
   U6143 : IVI port map( A => n2093, Z => n8245);
   U6144 : IVI port map( A => n1936, Z => n8246);
   U6145 : IVI port map( A => n1934, Z => n8247);
   U6146 : IVI port map( A => n2036, Z => n8248);
   U6147 : IVI port map( A => n2007, Z => n8249);
   U6148 : IVI port map( A => n2134, Z => n8250);
   U6149 : IVI port map( A => n2115, Z => n8253);
   U6150 : IVI port map( A => n2096, Z => n8254);
   U6151 : IVI port map( A => n1968, Z => n8255);
   U6152 : IVI port map( A => n1881, Z => n8256);
   U6153 : IVI port map( A => n2060, Z => n8258);
   U6154 : IVI port map( A => n2279, Z => n8261);
   U6155 : IVI port map( A => n2162, Z => n8266);
   U6156 : IVI port map( A => n2046, Z => n8268);
   U6157 : IVI port map( A => n2056, Z => n8269);
   U6158 : IVI port map( A => n1990, Z => n8270);
   U6159 : IVI port map( A => n1867, Z => n8271);
   U6160 : IVI port map( A => n2013, Z => n8272);
   U6161 : IVI port map( A => n1925, Z => n8273);
   U6162 : IVI port map( A => n1894, Z => n8274);
   U6163 : IVI port map( A => n149, Z => n8275);
   U6164 : IVI port map( A => n154, Z => n8276);
   U6165 : IVI port map( A => n108, Z => n8277);
   U6166 : IVI port map( A => n113, Z => n8278);
   U6167 : IVI port map( A => n172, Z => n8279);
   U6168 : IVI port map( A => n259, Z => n8280);
   U6169 : IVI port map( A => n58, Z => n8281);
   U6170 : IVI port map( A => n2281, Z => n8282);
   U6171 : IVI port map( A => n293, Z => n8283);
   U6172 : IVI port map( A => n286, Z => n8284);
   U6173 : IVI port map( A => n2476, Z => n8285);
   U6174 : IVI port map( A => n155, Z => n8286);
   U6175 : IVI port map( A => n280, Z => n8287);
   U6176 : IVI port map( A => n2033, Z => n8288);
   U6177 : IVI port map( A => n2278, Z => n8289);
   U6178 : IVI port map( A => n257, Z => n8290);
   U6179 : IVI port map( A => n1843, Z => n8291);
   U6180 : IVI port map( A => n1844, Z => n8292);
   U6181 : IVI port map( A => n1833, Z => n8293);
   U6182 : IVI port map( A => n1834, Z => n8294);
   U6183 : IVI port map( A => n1805, Z => n8295);
   U6184 : IVI port map( A => n1806, Z => n8296);
   U6185 : IVI port map( A => n2467, Z => n8297);
   U6186 : IVI port map( A => VALID_KEY_I, Z => n8298);
   U6187 : IVI port map( A => n336, Z => n8299);
   U6188 : IVI port map( A => RESET_I, Z => n8300);
   U6189 : IVI port map( A => n2483, Z => n8301);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_aes_dec_KEY_SIZE2.all;

entity aes_dec_KEY_SIZE2 is

   port( DATA_I : in std_logic_vector (7 downto 0);  VALID_DATA_I : in 
         std_logic;  KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, 
         RESET_I, CLK_I, CE_I : in std_logic;  KEY_READY_O, VALID_O : out 
         std_logic;  DATA_O : out std_logic_vector (7 downto 0));

end aes_dec_KEY_SIZE2;

architecture SYN_Behavioral of aes_dec_KEY_SIZE2 is

   component IVI
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EO
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EN
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO7
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component IV
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EON1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component IVDA
      port( A : in std_logic;  Y, Z : out std_logic);
   end component;
   
   component AO3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component NR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EOI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component EO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component ENI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2P
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4P
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component NR3P
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component key_expansion
      port( KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, CLK_I, 
            RESET_I, CE_I : in std_logic;  DONE_O : out std_logic;  GET_KEY_I :
            in std_logic;  KEY_NUMB_I : in std_logic_vector (5 downto 0);  
            KEY_EXP_O : out std_logic_vector (31 downto 0));
   end component;
   
   component NR4P
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO1P
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FD1
      port( D, CP : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_O_7_port, DATA_O_6_port, DATA_O_5_port, DATA_O_4_port, 
      DATA_O_3_port, DATA_O_2_port, DATA_O_1_port, DATA_O_0_port, GET_KEY, 
      v_INV_KEY_NUMB_5_port, v_INV_KEY_NUMB_4_port, v_INV_KEY_NUMB_3_port, 
      v_INV_KEY_NUMB_2_port, v_KEY_COLUMN_31_port, v_KEY_COLUMN_30_port, 
      v_KEY_COLUMN_29_port, v_KEY_COLUMN_28_port, v_KEY_COLUMN_27_port, 
      v_KEY_COLUMN_26_port, v_KEY_COLUMN_25_port, v_KEY_COLUMN_24_port, 
      v_KEY_COLUMN_23_port, v_KEY_COLUMN_22_port, v_KEY_COLUMN_21_port, 
      v_KEY_COLUMN_20_port, v_KEY_COLUMN_19_port, v_KEY_COLUMN_18_port, 
      v_KEY_COLUMN_17_port, v_KEY_COLUMN_16_port, v_KEY_COLUMN_15_port, 
      v_KEY_COLUMN_14_port, v_KEY_COLUMN_13_port, v_KEY_COLUMN_12_port, 
      v_KEY_COLUMN_11_port, v_KEY_COLUMN_10_port, v_KEY_COLUMN_9_port, 
      v_KEY_COLUMN_8_port, v_KEY_COLUMN_7_port, v_KEY_COLUMN_6_port, 
      v_KEY_COLUMN_5_port, v_KEY_COLUMN_4_port, v_KEY_COLUMN_3_port, 
      v_KEY_COLUMN_2_port, v_KEY_COLUMN_1_port, v_KEY_COLUMN_0_port, 
      v_CNT4_1_port, v_CNT4_0_port, v_DATA_COLUMN_31_port, 
      v_DATA_COLUMN_30_port, v_DATA_COLUMN_29_port, v_DATA_COLUMN_28_port, 
      v_DATA_COLUMN_27_port, v_DATA_COLUMN_26_port, v_DATA_COLUMN_25_port, 
      v_DATA_COLUMN_24_port, v_DATA_COLUMN_23_port, v_DATA_COLUMN_22_port, 
      v_DATA_COLUMN_21_port, v_DATA_COLUMN_20_port, v_DATA_COLUMN_19_port, 
      v_DATA_COLUMN_18_port, v_DATA_COLUMN_17_port, v_DATA_COLUMN_15_port, 
      v_DATA_COLUMN_14_port, v_DATA_COLUMN_13_port, v_DATA_COLUMN_12_port, 
      v_DATA_COLUMN_11_port, v_DATA_COLUMN_10_port, v_DATA_COLUMN_9_port, 
      v_DATA_COLUMN_7_port, v_DATA_COLUMN_6_port, v_DATA_COLUMN_5_port, 
      v_DATA_COLUMN_4_port, v_DATA_COLUMN_3_port, v_DATA_COLUMN_2_port, 
      v_DATA_COLUMN_1_port, v_CALCULATION_CNTR_7_port, 
      v_CALCULATION_CNTR_6_port, v_CALCULATION_CNTR_5_port, 
      v_CALCULATION_CNTR_4_port, v_CALCULATION_CNTR_3_port, 
      v_CALCULATION_CNTR_2_port, v_CALCULATION_CNTR_1_port, 
      v_CALCULATION_CNTR_0_port, N192, N199, N200, N201, N202, N203, 
      t_STATE_RAM0_0_31_port, t_STATE_RAM0_0_30_port, t_STATE_RAM0_0_29_port, 
      t_STATE_RAM0_0_28_port, t_STATE_RAM0_0_27_port, t_STATE_RAM0_0_26_port, 
      t_STATE_RAM0_0_25_port, t_STATE_RAM0_0_24_port, t_STATE_RAM0_0_23_port, 
      t_STATE_RAM0_0_22_port, t_STATE_RAM0_0_21_port, t_STATE_RAM0_0_20_port, 
      t_STATE_RAM0_0_19_port, t_STATE_RAM0_0_18_port, t_STATE_RAM0_0_17_port, 
      t_STATE_RAM0_0_16_port, t_STATE_RAM0_0_15_port, t_STATE_RAM0_0_14_port, 
      t_STATE_RAM0_0_13_port, t_STATE_RAM0_0_12_port, t_STATE_RAM0_0_11_port, 
      t_STATE_RAM0_0_10_port, t_STATE_RAM0_0_9_port, t_STATE_RAM0_0_8_port, 
      t_STATE_RAM0_0_7_port, t_STATE_RAM0_0_6_port, t_STATE_RAM0_0_5_port, 
      t_STATE_RAM0_0_4_port, t_STATE_RAM0_0_3_port, t_STATE_RAM0_0_2_port, 
      t_STATE_RAM0_0_1_port, t_STATE_RAM0_0_0_port, t_STATE_RAM0_1_31_port, 
      t_STATE_RAM0_1_30_port, t_STATE_RAM0_1_29_port, t_STATE_RAM0_1_28_port, 
      t_STATE_RAM0_1_27_port, t_STATE_RAM0_1_26_port, t_STATE_RAM0_1_25_port, 
      t_STATE_RAM0_1_24_port, t_STATE_RAM0_1_23_port, t_STATE_RAM0_1_22_port, 
      t_STATE_RAM0_1_21_port, t_STATE_RAM0_1_20_port, t_STATE_RAM0_1_19_port, 
      t_STATE_RAM0_1_18_port, t_STATE_RAM0_1_17_port, t_STATE_RAM0_1_16_port, 
      t_STATE_RAM0_1_15_port, t_STATE_RAM0_1_14_port, t_STATE_RAM0_1_13_port, 
      t_STATE_RAM0_1_12_port, t_STATE_RAM0_1_11_port, t_STATE_RAM0_1_10_port, 
      t_STATE_RAM0_1_9_port, t_STATE_RAM0_1_8_port, t_STATE_RAM0_1_7_port, 
      t_STATE_RAM0_1_6_port, t_STATE_RAM0_1_5_port, t_STATE_RAM0_1_4_port, 
      t_STATE_RAM0_1_3_port, t_STATE_RAM0_1_2_port, t_STATE_RAM0_1_1_port, 
      t_STATE_RAM0_1_0_port, t_STATE_RAM0_2_31_port, t_STATE_RAM0_2_30_port, 
      t_STATE_RAM0_2_29_port, t_STATE_RAM0_2_28_port, t_STATE_RAM0_2_27_port, 
      t_STATE_RAM0_2_26_port, t_STATE_RAM0_2_25_port, t_STATE_RAM0_2_24_port, 
      t_STATE_RAM0_2_23_port, t_STATE_RAM0_2_22_port, t_STATE_RAM0_2_21_port, 
      t_STATE_RAM0_2_20_port, t_STATE_RAM0_2_19_port, t_STATE_RAM0_2_18_port, 
      t_STATE_RAM0_2_17_port, t_STATE_RAM0_2_16_port, t_STATE_RAM0_2_15_port, 
      t_STATE_RAM0_2_14_port, t_STATE_RAM0_2_13_port, t_STATE_RAM0_2_12_port, 
      t_STATE_RAM0_2_11_port, t_STATE_RAM0_2_10_port, t_STATE_RAM0_2_9_port, 
      t_STATE_RAM0_2_8_port, t_STATE_RAM0_2_7_port, t_STATE_RAM0_2_6_port, 
      t_STATE_RAM0_2_5_port, t_STATE_RAM0_2_4_port, t_STATE_RAM0_2_3_port, 
      t_STATE_RAM0_2_2_port, t_STATE_RAM0_2_1_port, t_STATE_RAM0_2_0_port, 
      v_RAM_OUT0_31_port, v_RAM_OUT0_30_port, v_RAM_OUT0_29_port, 
      v_RAM_OUT0_28_port, v_RAM_OUT0_27_port, v_RAM_OUT0_26_port, 
      v_RAM_OUT0_25_port, v_RAM_OUT0_24_port, v_RAM_OUT0_23_port, 
      v_RAM_OUT0_22_port, v_RAM_OUT0_21_port, v_RAM_OUT0_20_port, 
      v_RAM_OUT0_19_port, v_RAM_OUT0_18_port, v_RAM_OUT0_17_port, 
      v_RAM_OUT0_16_port, v_RAM_OUT0_15_port, v_RAM_OUT0_14_port, 
      v_RAM_OUT0_13_port, v_RAM_OUT0_12_port, v_RAM_OUT0_11_port, 
      v_RAM_OUT0_10_port, v_RAM_OUT0_9_port, v_RAM_OUT0_7_port, 
      v_RAM_OUT0_6_port, v_RAM_OUT0_5_port, v_RAM_OUT0_4_port, 
      v_RAM_OUT0_3_port, v_RAM_OUT0_2_port, v_RAM_OUT0_1_port, 
      v_RAM_OUT0_0_port, N2083, N2084, N2085, N2086, N2087, N2088, N2089, n3, 
      n4, n10, n11, n13, n14, n16, n17, n19, n20, n22, n23, n25, n26, n28, n29,
      n31, n32, n34, n35, n37, n38, n40, n41, n43, n44, n46, n47, n49, n50, n52
      , n53, n55, n56, n58, n59, n61, n62, n64, n65, n67, n68, n70, n71, n73, 
      n74, n76, n77, n79, n80, n82, n83, n85, n86, n88, n89, n91, n92, n94, n95
      , n97, n98, n100, n101, n103, n105, n107, n108, n109, n111, n113, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n135, n136, n138, n139, n140, n141, 
      n142, n143, n145, n146, n147, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n188, n189, n190, n191, n192_port, 
      n193, n196, n197, n198, n199_port, n200_port, n201_port, n204, n205, n206
      , n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, 
      n417, n418, n419, n420, n421, n423, n424, n425, n426, n427, n428, n429, 
      n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n555, n556, n557, n558, n559, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n611, n612, n613, n614, n615, n616, n618, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, 
      n659, n660, n661, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n691, n692, n694, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n725, n726, n727, n728, n729, n730, n731, n732, n733, n735, n736, 
      n737, n738, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
      n750, n751, n752, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n828, n829, n830, n831, n832, n834, n835, n836, n837, n838, 
      n839, n840, n841, n842, n843, n844, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, 
      n878, n879, n881, n882, n883, n884, n885, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n941, 
      n942, n943, n944, n945, n946, n947, n949, n950, n951, n952, n953, n954, 
      n955, n957, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, 
      n982, n983, n984, n985, n986, n987, n988, n989, n991, n992, n993, n994, 
      n995, n996, n998, n999, n1000, n1001, n1002, n1003, n1005, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1019, n1020, n1021, 
      n1022, n1026, n1027, n1028, n1029, n1031, n1032, n1033, n1034, n1035, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1048, 
      n1049, n1050, n1051, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1078, n1079, n1080, n1081, n1082, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1114, n1115, n1116, n1117, n1118, n1121, 
      n1122, n1123, n1124, n1127, n1128, n1129, n1130, n1131, n1133, n1134, 
      n1135, n1136, n1139, n1140, n1141, n1142, n1143, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1152, n1153, n1154, n1155, n1156, n1160, n1161, 
      n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1171, n1172, n1174, 
      n1175, n1178, n1179, n1180, n1183, n1184, n1185, n1186, n1188, n1189, 
      n1191, n1194, n1195, n1196, n1197, n1200, n1201, n1202, n1203, n1206, 
      n1209, n1210, n1212, n1213, n1216, n1217, n1218, n1219, n1221, n1222, 
      n1223, n1227, n1228, n1229, n1231, n1232, n1237, n1238, n1241, n1242, 
      n1243, n1245, n1246, n1250, n1251, n1254, n1255, n1256, n1258, n1259, 
      n1263, n1264, n1265, n1266, n1268, n1269, n1270, n1271, n1272, n1273, 
      n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1301, n1302, 
      n1303, n1304, n1305, n1315, n1319, n1320, n1330, n1331, n1332, n1333, 
      n1335, n1336, n1339, n1340, n1342, n1343, n1348, n1349, n1353, n1354, 
      n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1365, n1366, 
      n1369, n1370, n1372, n1373, n1374, n1375, n1376, n1377, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1406, n1407, n1409, n1410, n1411, n1413, n1418, 
      n1424, n1426, n1428, n1429, n1430, n1433, n1434, n1435, n1436, n1439, 
      n1440, n1441, n1444, n1445, n1446, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1457, n1458, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1469, n1470, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1491, n1492, n1493, n1494, n1497, n1498, n1499, n1500, 
      n1501, n1502, n1503, n1504, n1506, n1507, n1508, n1509, n1511, n1512, 
      n1513, n1514, n1516, n1517, n1518, n1519, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1529, n1530, n1531, n1532, n1533, n1534, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1544, n1545, n1546, n1547, n1550, n1551, 
      n1552, n1553, n1556, n1557, n1558, n1559, n1561, n1562, n1563, n1564, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1579, n1581, n1582, n1583, n1584, n1585, n1586, n1589, 
      n1590, n1591, n1592, n1594, n1595, n1596, n1597, n1600, n1601, n1602, 
      n1603, n1605, n1606, n1607, n1608, n1610, n1611, n1612, n1613, n1614, 
      n1616, n1617, n1618, n1619, n1620, n1622, n1624, n1625, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1637, n1638, n1639, n1640, 
      n1641, n1644, n1648, n1649, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1663, n1664, n1665, n1667, n1668, n1669, n1670, n1671, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1682, n1683, n1684, n1685, n1688, n1689, 
      n1691, n1692, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, 
      n1702, n1703, n1704, n1705, n1706, n1707, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
      n1734, n1735, n1736, n1737, n1738, n1739, n1741, n1742, n1743, n1745, 
      n1746, n1747, n1749, n1750, n1751, n1753, n1754, n1755, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1772, n1773, n1774, n1775, n1776, n1777, n1779, n1780, 
      n1781, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, 
      n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
      n1802, n1804, n1805, n1806, n1807, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
      n1825, n1826, n1827, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1841, n1843, n1844, n1845, n1848, n1852, 
      n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1862, n1863, n1864, 
      n1865, n1866, n1868, n1869, n1873, n1874, n1875, n1876, n1878, n1879, 
      n1880, n1881, n1882, n1884, n1887, n1888, n1889, n1890, n1892, n1893, 
      n1894, n1895, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n1905, n1906, n1908, n1909, n1910, n1911, n1912, n1913, n1915, n1917, 
      n1919, n1920, n1922, n1923, n1924, n1926, n1927, n1928, n1929, n1930, 
      n1931, n1933, n1935, n1936, n1938, n1939, n1940, n1941, n1942, n1943, 
      n1944, n1945, n1946, n1949, n1950, n1951, n1953, n1954, n1956, n1958, 
      n1959, n1961, n1962, n1963, n1964, n1966, n1967, n1968, n1969, n1971, 
      n1972, n1974, n1976, n1978, n1979, n1980, n1981, n1982, n1984, n1985, 
      n1986, n1988, n1989, n1990, n1992, n1993, n1994, n1995, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2012, n2015, n2018, n2021, n2023, n2026, n2027, n2028, 
      n2029, n2030, n2032, n2033, n2034, n2035, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2046, n2047, n2049, n2050, n2051, n2053, n2054, n2055, 
      n2056, n2057, n2059, n2060, n2062, n2063, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2075, n2076, n2077, n2078, n2079, 
      n2080, n2081, n2082, n2083_port, n2084_port, n2085_port, n2086_port, 
      n2088_port, n2089_port, n2090, n2091, n2092, n2093, n2094, n2095, n2097, 
      n2098, n2101, n2102, n2108, n2109, n2110, n2111, n2112, n2113, n2114, 
      n2116, n2117, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2138, 
      n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
      n2149, n2150, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2160, 
      n2161, n2162, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, 
      n2172, n2173, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
      n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, 
      n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2222, n2223, n2224, n2225, 
      n2227, n2228, n2229, n2230, n2231, n2233, n2234, n2235, n2236, n2238, 
      n2239, n2240, n2241, n2242, n2243, n2244, n2246, n2248, n2249, n2250, 
      n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, 
      n2261, n2262, n2263, n2264, n2265, n2267, n2268, n2269, n2270, n2271, 
      n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2298, n2301, n2302, n2303, n2304, n2305, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2332, n2334, n2335, n2336, n2337, n2338, 
      n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, 
      n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, 
      n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
      n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, 
      n2380, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2390, n2391, 
      n2392, n2393, n2394, n2395, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2419, n2420, n2421, n2423, n2424, 
      n2425, n2427, n2428, n2429, n2430, n2431, n2433, n2437, n2438, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2452, n2453, n2455, n2456, n2457, 
      n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2467, n2468, n2469, 
      n2470, n2473, n2474, n2476, n2477, n2479, n2480, n2481, n2482, n2483, 
      n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, 
      n2494, n2495, n2497, n2499, n2501, n2502, n2505, n2507, n2508, n2509, 
      n2511, n2512, n2513, n2515, n2516, n2517, n2519, n2520, n2521, n2522, 
      n2524, n2525, n2526, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2536, n2539, n2540, n2541, n2542, n2544, n2545, n2546, n2547, n2549, 
      n2550, n2551, n2552, n2553, n2556, n2558, n2559, n2561, n2562, n2563, 
      n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
      n2574, n2575, n2577, n2578, n2579, n2581, n2582, n2583, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2592, n2593, n2597, n2598, n2600, n2601, 
      n2602, n2604, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, 
      n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2625, 
      n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, 
      n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2657, 
      n2658, n2659, n2662, n2664, n2665, n2666, n2667, n2668, n2669, n2670, 
      n2671, n2672, n2674, n2675, n2676, n2677, n2679, n2680, n2681, n2682, 
      n2683, n2684, n2685, n2686, n2689, n2690, n2692, n2693, n2694, n2695, 
      n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2706, 
      n2707, n2708, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
      n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2769, n2770, 
      n2771, n2772, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, 
      n2782, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
      n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, 
      n2803, n2804, n2805, n2806, n2807, n2808, n2810, n2811, n2812, n2813, 
      n2814, n2815, n2817, n2818, n2820, n2821, n2822, n2823, n2824, n2825, 
      n2826, n2827, n2828, n2829, n2830, n2832, n2833, n2835, n2836, n2837, 
      n2838, n2839, n2840, n2841, n2842, n2843, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2871, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
      n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, 
      n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
      n2901, n2902, n2903, n2905, n2906, n2908, n2909, n2912, n2914, n2915, 
      n2916, n2918, n2919, n2920, n2922, n2924, n2925, n2927, n2928, n2930, 
      n2931, n2932, n2934, n2935, n2936, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2945, n2947, n2948, n2949, n2950, n2951, n2952, n2954, n2955, 
      n2957, n2958, n2959, n2960, n2961, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2976, n2977, n2978, n2979, 
      n2980, n2981, n2982, n2984, n2985, n2986, n2988, n2989, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2998, n2999, n3003, n3004, n3005, n3007, 
      n3008, n3009, n3010, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
      n3020, n3021, n3022, n3023, n3024, n3026, n3027, n3028, n3029, n3030, 
      n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, 
      n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3051, n3052, 
      n3053, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3065, n3066, n3067, n3070, n3072, n3073, n3074, n3075, n3076, n3077, 
      n3078, n3079, n3080, n3082, n3083, n3084, n3085, n3087, n3088, n3089, 
      n3090, n3091, n3092, n3093, n3094, n3097, n3098, n3099, n3100, n3101, 
      n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
      n3112, n3113, n3114, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, 
      n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, 
      n3165, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3176, 
      n3177, n3178, n3179, n3181, n3182, n3183, n3184, n3185, n3186, n3187, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3206, n3207, n3208, n3209, 
      n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3218, n3219, n3220, 
      n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
      n3231, n3232, n3233, n3234, n3235, n3237, n3238, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
      n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, 
      n3274, n3275, n3276, n3277, n3278, n3279, n3281, n3282, n3283, n3284, 
      n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
      n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, 
      n3305, n3306, n3308, n3309, n3310, n3311, n3312, n3315, n3317, n3318, 
      n3319, n3321, n3322, n3323, n3325, n3327, n3328, n3330, n3331, n3333, 
      n3334, n3335, n3337, n3338, n3339, n3341, n3342, n3343, n3344, n3345, 
      n3346, n3348, n3350, n3351, n3352, n3353, n3354, n3355, n3357, n3358, 
      n3360, n3361, n3362, n3363, n3364, n3367, n3368, n3369, n3370, n3371, 
      n3372, n3373, n3374, n3375, n3376, n3377, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3387, n3388, n3389, n3391, n3392, n3394, n3395, 
      n3396, n3397, n3398, n3399, n3401, n3402, n3406, n3407, n3408, n3410, 
      n3411, n3412, n3413, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3429, n3430, n3431, n3432, n3433, 
      n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, 
      n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3454, n3455, 
      n3456, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3468, n3469, n3470, n3473, n3475, n3476, n3477, n3478, n3479, n3480, 
      n3481, n3482, n3483, n3485, n3486, n3487, n3488, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3500, n3501, n3503, n3504, n3505, 
      n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, 
      n3516, n3517, n3518, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3537, 
      n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3580, 
      n3581, n3582, n3583, n3585, n3586, n3587, n3588, n3589, n3590, n3591, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3610, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3622, n3623, n3624, 
      n3625, n3626, n3627, n3628, n3630, n3631, n3632, n3633, n3634, n3635, 
      n3636, n3637, n3638, n3639, n3640, n3642, n3643, n3645, n3646, n3647, 
      n3648, n3649, n3650, n3651, n3652, n3653, n3655, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, 
      n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3689, n3690, 
      n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, 
      n3701, n3703, n3704, n3705, n3706, n3708, n3710, n3712, n3713, n3714, 
      n3715, n3716, n3717, n3720, n3721, n3722, n3723, n3724, n3725, n3726, 
      n3727, n3728, n3729, n3730, n3731, n3733, n3734, n3735, n3736, n3737, 
      n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, 
      n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, 
      n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, 
      n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, 
      n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3809, n3810, 
      n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, 
      n3821, n3823, n3824, n3825, n3827, n3828, n3829, n3835, n3838, n3839, 
      n3840, n3841, n3842, n3843, n3844, n3845, n3847, n3848, n3850, n3854, 
      n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3867, 
      n3870, n3871, n3872, n3873, n3874, n3879, n3880, n3882, n3886, n3888, 
      n3889, n3894, n3899, n3902, n3903, n3904, n3905, n3906, n3907, n3908, 
      n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
      n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3931, 
      n3934, n3935, n3936, n3937, n3938, n3942, n3943, n3944, n3945, n3946, 
      n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, 
      n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
      n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, 
      n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, 
      n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, 
      n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, 
      n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, 
      n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, 
      n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, 
      n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
      n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, 
      n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
      n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, 
      n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, 
      n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
      n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, 
      n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, 
      n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
      n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, 
      n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
      n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, 
      n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, 
      n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, 
      n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
      n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, 
      n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, 
      n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, 
      n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
      n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, 
      n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, 
      n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
      n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
      n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, 
      n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, 
      n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
      n4297, n4298, n4299, n4300, n4301, n4303, n4304, n4305, n4309, n4310, 
      n4311, n4312, n4313, n4314, n4315, n4323, n4331, n4339, n4340, n4348, 
      n4349, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, 
      n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, 
      n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, 
      n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, 
      n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, 
      n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, 
      n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, 
      n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, 
      n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
      n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, 
      n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, 
      n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, 
      n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, 
      n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, 
      n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, 
      n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, 
      n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, 
      n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, 
      n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, 
      n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, 
      n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, 
      n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, 
      n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, 
      n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, 
      n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, 
      n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, 
      n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, 
      n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, 
      n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, 
      n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
      n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, 
      n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, 
      n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, 
      n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, 
      n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, 
      n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, 
      n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, 
      n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, 
      n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, 
      n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, 
      n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, 
      n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, 
      n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, 
      n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, 
      n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, 
      n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, 
      n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, 
      n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, 
      n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, 
      n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, 
      n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, 
      n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, 
      n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, 
      n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, 
      n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, 
      n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, 
      n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, 
      n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, 
      n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, 
      n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, 
      n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, 
      n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, 
      n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, 
      n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, 
      n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, 
      n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, 
      n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, 
      n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, 
      n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, 
      n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, 
      n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, 
      n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, 
      n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, 
      n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, 
      n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, 
      n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, 
      n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, 
      n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, 
      n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, 
      n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, 
      n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, 
      n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, 
      n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, 
      n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, 
      n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, 
      n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, 
      n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, 
      n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, 
      n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, 
      n5241, n5242, n5243, n5244, n5245, n5246, n_3137, n_3138, n_3139, n_3140,
      n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, 
      n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, 
      n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, 
      n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, 
      n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, 
      n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, 
      n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, 
      n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, 
      n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, 
      n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, 
      n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, 
      n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, 
      n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, 
      n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, 
      n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, 
      n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, 
      n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, 
      n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, 
      n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, 
      n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, 
      n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, 
      n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, 
      n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, 
      n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, 
      n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, 
      n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, 
      n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, 
      n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, 
      n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, 
      n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, 
      n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, 
      n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, 
      n_3429, n_3430, n_3431 : std_logic;

begin
   DATA_O <= ( DATA_O_7_port, DATA_O_6_port, DATA_O_5_port, DATA_O_4_port, 
      DATA_O_3_port, DATA_O_2_port, DATA_O_1_port, DATA_O_0_port );
   
   GET_KEY_reg : FD1 port map( D => N192, CP => CLK_I, Q => GET_KEY, QN => 
                           n3952);
   v_CNT4_reg_0_inst : FD1 port map( D => n4349, CP => CLK_I, Q => 
                           v_CNT4_0_port, QN => n4380);
   v_DATA_COLUMN_reg_24_inst : FD1 port map( D => n4348, CP => CLK_I, Q => 
                           v_DATA_COLUMN_24_port, QN => n_3137);
   v_DATA_COLUMN_reg_25_inst : FD1 port map( D => n4995, CP => CLK_I, Q => 
                           v_DATA_COLUMN_25_port, QN => n_3138);
   v_DATA_COLUMN_reg_26_inst : FD1 port map( D => n4991, CP => CLK_I, Q => 
                           v_DATA_COLUMN_26_port, QN => n_3139);
   v_DATA_COLUMN_reg_27_inst : FD1 port map( D => n4987, CP => CLK_I, Q => 
                           v_DATA_COLUMN_27_port, QN => n_3140);
   v_DATA_COLUMN_reg_28_inst : FD1 port map( D => n4983, CP => CLK_I, Q => 
                           v_DATA_COLUMN_28_port, QN => n_3141);
   v_DATA_COLUMN_reg_29_inst : FD1 port map( D => n4979, CP => CLK_I, Q => 
                           v_DATA_COLUMN_29_port, QN => n_3142);
   v_DATA_COLUMN_reg_30_inst : FD1 port map( D => n4975, CP => CLK_I, Q => 
                           v_DATA_COLUMN_30_port, QN => n_3143);
   v_DATA_COLUMN_reg_31_inst : FD1 port map( D => n4971, CP => CLK_I, Q => 
                           v_DATA_COLUMN_31_port, QN => n_3144);
   v_CNT4_reg_1_inst : FD1 port map( D => n4340, CP => CLK_I, Q => 
                           v_CNT4_1_port, QN => n4540);
   v_DATA_COLUMN_reg_8_inst : FD1 port map( D => n4339, CP => CLK_I, Q => 
                           n_3145, QN => n4602);
   v_DATA_COLUMN_reg_9_inst : FD1 port map( D => n4994, CP => CLK_I, Q => 
                           v_DATA_COLUMN_9_port, QN => n_3146);
   v_DATA_COLUMN_reg_10_inst : FD1 port map( D => n4993, CP => CLK_I, Q => 
                           v_DATA_COLUMN_10_port, QN => n_3147);
   v_DATA_COLUMN_reg_11_inst : FD1 port map( D => n4989, CP => CLK_I, Q => 
                           v_DATA_COLUMN_11_port, QN => n_3148);
   v_DATA_COLUMN_reg_12_inst : FD1 port map( D => n4985, CP => CLK_I, Q => 
                           v_DATA_COLUMN_12_port, QN => n_3149);
   v_DATA_COLUMN_reg_13_inst : FD1 port map( D => n4981, CP => CLK_I, Q => 
                           v_DATA_COLUMN_13_port, QN => n_3150);
   v_DATA_COLUMN_reg_14_inst : FD1 port map( D => n4977, CP => CLK_I, Q => 
                           v_DATA_COLUMN_14_port, QN => n_3151);
   v_DATA_COLUMN_reg_15_inst : FD1 port map( D => n4973, CP => CLK_I, Q => 
                           v_DATA_COLUMN_15_port, QN => n_3152);
   v_DATA_COLUMN_reg_16_inst : FD1 port map( D => n4331, CP => CLK_I, Q => 
                           n_3153, QN => n4601);
   v_DATA_COLUMN_reg_17_inst : FD1 port map( D => n4997, CP => CLK_I, Q => 
                           v_DATA_COLUMN_17_port, QN => n_3154);
   v_DATA_COLUMN_reg_18_inst : FD1 port map( D => n4992, CP => CLK_I, Q => 
                           v_DATA_COLUMN_18_port, QN => n_3155);
   v_DATA_COLUMN_reg_19_inst : FD1 port map( D => n4988, CP => CLK_I, Q => 
                           v_DATA_COLUMN_19_port, QN => n_3156);
   v_DATA_COLUMN_reg_20_inst : FD1 port map( D => n4984, CP => CLK_I, Q => 
                           v_DATA_COLUMN_20_port, QN => n_3157);
   v_DATA_COLUMN_reg_21_inst : FD1 port map( D => n4980, CP => CLK_I, Q => 
                           v_DATA_COLUMN_21_port, QN => n_3158);
   v_DATA_COLUMN_reg_22_inst : FD1 port map( D => n4976, CP => CLK_I, Q => 
                           v_DATA_COLUMN_22_port, QN => n_3159);
   v_DATA_COLUMN_reg_23_inst : FD1 port map( D => n4972, CP => CLK_I, Q => 
                           v_DATA_COLUMN_23_port, QN => n_3160);
   v_DATA_COLUMN_reg_0_inst : FD1 port map( D => n4323, CP => CLK_I, Q => 
                           n_3161, QN => n4600);
   v_DATA_COLUMN_reg_1_inst : FD1 port map( D => n4996, CP => CLK_I, Q => 
                           v_DATA_COLUMN_1_port, QN => n_3162);
   v_DATA_COLUMN_reg_2_inst : FD1 port map( D => n4990, CP => CLK_I, Q => 
                           v_DATA_COLUMN_2_port, QN => n_3163);
   v_DATA_COLUMN_reg_3_inst : FD1 port map( D => n4986, CP => CLK_I, Q => 
                           v_DATA_COLUMN_3_port, QN => n_3164);
   v_DATA_COLUMN_reg_4_inst : FD1 port map( D => n4982, CP => CLK_I, Q => 
                           v_DATA_COLUMN_4_port, QN => n_3165);
   v_DATA_COLUMN_reg_5_inst : FD1 port map( D => n4978, CP => CLK_I, Q => 
                           v_DATA_COLUMN_5_port, QN => n_3166);
   v_DATA_COLUMN_reg_6_inst : FD1 port map( D => n4974, CP => CLK_I, Q => 
                           v_DATA_COLUMN_6_port, QN => n_3167);
   v_DATA_COLUMN_reg_7_inst : FD1 port map( D => n4970, CP => CLK_I, Q => 
                           v_DATA_COLUMN_7_port, QN => n_3168);
   FF_VALID_DATA_reg : FD1 port map( D => n4315, CP => CLK_I, Q => n4414, QN =>
                           n3959);
   LAST_ROUND_reg : FD1 port map( D => n4314, CP => CLK_I, Q => n4439, QN => 
                           n3958);
   v_CALCULATION_CNTR_reg_0_inst : FD1 port map( D => n4313, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_0_port, QN => n4604);
   v_CALCULATION_CNTR_reg_1_inst : FD1 port map( D => n4312, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_1_port, QN => n4411);
   v_CALCULATION_CNTR_reg_2_inst : FD1 port map( D => n4311, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_2_port, QN => n4556);
   v_CALCULATION_CNTR_reg_3_inst : FD1 port map( D => n4310, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_3_port, QN => n4369);
   v_CALCULATION_CNTR_reg_4_inst : FD1 port map( D => n4309, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_4_port, QN => n4527);
   v_CALCULATION_CNTR_reg_5_inst : FD1 port map( D => n5008, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_5_port, QN => n_3169);
   v_CALCULATION_CNTR_reg_6_inst : FD1 port map( D => n5007, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_6_port, QN => n4599);
   v_CALCULATION_CNTR_reg_7_inst : FD1 port map( D => n5006, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_7_port, QN => n_3170);
   FF_GET_KEY_reg : FD1 port map( D => n4305, CP => CLK_I, Q => n_3171, QN => 
                           n3951);
   SRAM_WREN0_reg : FD1 port map( D => n4304, CP => CLK_I, Q => n_3172, QN => 
                           n3950);
   i_RAM_ADDR_WR0_reg_0_inst : FD1 port map( D => n4303, CP => CLK_I, Q => 
                           n_3173, QN => n3949);
   i_RAM_ADDR_WR0_reg_1_inst : FD1 port map( D => n5001, CP => CLK_I, Q => 
                           n4466, QN => n3948);
   v_KEY_NUMB_reg_5_inst : FD1 port map( D => n4301, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_5_port, QN => n3947);
   v_KEY_NUMB_reg_0_inst : FD1 port map( D => n4300, CP => CLK_I, Q => n_3174, 
                           QN => n4667);
   v_KEY_NUMB_reg_1_inst : FD1 port map( D => n4299, CP => CLK_I, Q => n_3175, 
                           QN => n4666);
   v_KEY_NUMB_reg_2_inst : FD1 port map( D => n4298, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_2_port, QN => n3946);
   v_KEY_NUMB_reg_3_inst : FD1 port map( D => n4297, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_3_port, QN => n3945);
   v_KEY_NUMB_reg_4_inst : FD1 port map( D => n4296, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_4_port, QN => n3944);
   i_RAM_ADDR_RD0_reg_0_inst : FD1 port map( D => n4295, CP => CLK_I, Q => 
                           n4603, QN => n3943);
   i_RAM_ADDR_RD0_reg_1_inst : FD1 port map( D => n4294, CP => CLK_I, Q => 
                           n4366, QN => n3942);
   CALCULATION_reg : FD1 port map( D => n4293, CP => CLK_I, Q => n_3176, QN => 
                           n3957);
   i_ROUND_reg_0_inst : FD1 port map( D => n4292, CP => CLK_I, Q => n_3177, QN 
                           => n3954);
   i_ROUND_reg_1_inst : FD1 port map( D => n4291, CP => CLK_I, Q => n4471, QN 
                           => n3953);
   i_ROUND_reg_2_inst : FD1 port map( D => n4290, CP => CLK_I, Q => n4633, QN 
                           => n3955);
   i_ROUND_reg_3_inst : FD1 port map( D => n4289, CP => CLK_I, Q => n_3178, QN 
                           => n3956);
   STATE_TABLE1_reg_0_7_inst : FD1 port map( D => n4288, CP => CLK_I, Q => 
                           n4431, QN => n_3179);
   STATE_TABLE1_reg_0_6_inst : FD1 port map( D => n4287, CP => CLK_I, Q => 
                           n4406, QN => n_3180);
   STATE_TABLE1_reg_0_5_inst : FD1 port map( D => n4286, CP => CLK_I, Q => 
                           n4523, QN => n_3181);
   STATE_TABLE1_reg_0_4_inst : FD1 port map( D => n4285, CP => CLK_I, Q => 
                           n4609, QN => n3938);
   STATE_TABLE1_reg_0_3_inst : FD1 port map( D => n4284, CP => CLK_I, Q => 
                           n4608, QN => n3937);
   STATE_TABLE1_reg_0_2_inst : FD1 port map( D => n4283, CP => CLK_I, Q => 
                           n4607, QN => n3936);
   STATE_TABLE1_reg_0_1_inst : FD1 port map( D => n4282, CP => CLK_I, Q => 
                           n4606, QN => n3935);
   STATE_TABLE1_reg_0_0_inst : FD1 port map( D => n4281, CP => CLK_I, Q => 
                           n4605, QN => n3934);
   STATE_TABLE1_reg_1_7_inst : FD1 port map( D => n4280, CP => CLK_I, Q => 
                           n4407, QN => n_3182);
   STATE_TABLE1_reg_1_6_inst : FD1 port map( D => n4279, CP => CLK_I, Q => 
                           n4419, QN => n_3183);
   STATE_TABLE1_reg_1_5_inst : FD1 port map( D => n4278, CP => CLK_I, Q => 
                           n4612, QN => n3931);
   STATE_TABLE1_reg_1_4_inst : FD1 port map( D => n4277, CP => CLK_I, Q => 
                           n4551, QN => n_3184);
   STATE_TABLE1_reg_1_3_inst : FD1 port map( D => n4276, CP => CLK_I, Q => 
                           n4442, QN => n_3185);
   STATE_TABLE1_reg_1_2_inst : FD1 port map( D => n4275, CP => CLK_I, Q => 
                           n4418, QN => n_3186);
   STATE_TABLE1_reg_1_1_inst : FD1 port map( D => n4274, CP => CLK_I, Q => 
                           n4611, QN => n3927);
   STATE_TABLE1_reg_1_0_inst : FD1 port map( D => n4273, CP => CLK_I, Q => 
                           n4610, QN => n3926);
   STATE_TABLE1_reg_2_7_inst : FD1 port map( D => n4272, CP => CLK_I, Q => 
                           n4536, QN => n3925);
   STATE_TABLE1_reg_2_6_inst : FD1 port map( D => n4271, CP => CLK_I, Q => 
                           n4426, QN => n3924);
   STATE_TABLE1_reg_2_5_inst : FD1 port map( D => n4270, CP => CLK_I, Q => 
                           n4425, QN => n3923);
   STATE_TABLE1_reg_2_4_inst : FD1 port map( D => n4269, CP => CLK_I, Q => 
                           n4555, QN => n3922);
   STATE_TABLE1_reg_2_3_inst : FD1 port map( D => n4268, CP => CLK_I, Q => 
                           n4624, QN => n3921);
   STATE_TABLE1_reg_2_2_inst : FD1 port map( D => n4267, CP => CLK_I, Q => 
                           n4623, QN => n3920);
   STATE_TABLE1_reg_2_1_inst : FD1 port map( D => n4266, CP => CLK_I, Q => 
                           n4562, QN => n3919);
   STATE_TABLE1_reg_2_0_inst : FD1 port map( D => n4265, CP => CLK_I, Q => 
                           n4622, QN => n3918);
   STATE_TABLE1_reg_3_7_inst : FD1 port map( D => n4264, CP => CLK_I, Q => 
                           n4538, QN => n3917);
   STATE_TABLE1_reg_3_6_inst : FD1 port map( D => n4263, CP => CLK_I, Q => 
                           n4427, QN => n3916);
   STATE_TABLE1_reg_3_5_inst : FD1 port map( D => n4262, CP => CLK_I, Q => 
                           n4537, QN => n3915);
   STATE_TABLE1_reg_3_4_inst : FD1 port map( D => n4261, CP => CLK_I, Q => 
                           n4627, QN => n3914);
   STATE_TABLE1_reg_3_3_inst : FD1 port map( D => n4260, CP => CLK_I, Q => 
                           n4449, QN => n3913);
   STATE_TABLE1_reg_3_2_inst : FD1 port map( D => n4259, CP => CLK_I, Q => 
                           n4626, QN => n3912);
   STATE_TABLE1_reg_3_1_inst : FD1 port map( D => n4258, CP => CLK_I, Q => 
                           n4625, QN => n3911);
   STATE_TABLE1_reg_3_0_inst : FD1 port map( D => n4257, CP => CLK_I, Q => 
                           n4440, QN => n3910);
   STATE_TABLE1_reg_4_7_inst : FD1 port map( D => n4256, CP => CLK_I, Q => 
                           n4450, QN => n3909);
   STATE_TABLE1_reg_4_6_inst : FD1 port map( D => n4255, CP => CLK_I, Q => 
                           n4539, QN => n3908);
   STATE_TABLE1_reg_4_5_inst : FD1 port map( D => n4254, CP => CLK_I, Q => 
                           n4526, QN => n3907);
   STATE_TABLE1_reg_4_4_inst : FD1 port map( D => n4253, CP => CLK_I, Q => 
                           n4632, QN => n3906);
   STATE_TABLE1_reg_4_3_inst : FD1 port map( D => n4252, CP => CLK_I, Q => 
                           n4631, QN => n3905);
   STATE_TABLE1_reg_4_2_inst : FD1 port map( D => n4251, CP => CLK_I, Q => 
                           n4630, QN => n3904);
   STATE_TABLE1_reg_4_1_inst : FD1 port map( D => n4250, CP => CLK_I, Q => 
                           n4629, QN => n3903);
   STATE_TABLE1_reg_4_0_inst : FD1 port map( D => n4249, CP => CLK_I, Q => 
                           n4628, QN => n3902);
   STATE_TABLE1_reg_5_7_inst : FD1 port map( D => n4248, CP => CLK_I, Q => 
                           n4420, QN => n_3187);
   STATE_TABLE1_reg_5_6_inst : FD1 port map( D => n4247, CP => CLK_I, Q => 
                           n4384, QN => n_3188);
   STATE_TABLE1_reg_5_5_inst : FD1 port map( D => n4246, CP => CLK_I, Q => 
                           n4572, QN => n3899);
   STATE_TABLE1_reg_5_4_inst : FD1 port map( D => n4245, CP => CLK_I, Q => 
                           n4453, QN => n_3189);
   STATE_TABLE1_reg_5_3_inst : FD1 port map( D => n4244, CP => CLK_I, Q => 
                           n4452, QN => n_3190);
   STATE_TABLE1_reg_5_2_inst : FD1 port map( D => n4243, CP => CLK_I, Q => 
                           n4436, QN => n_3191);
   STATE_TABLE1_reg_5_1_inst : FD1 port map( D => n4242, CP => CLK_I, Q => 
                           n4443, QN => n_3192);
   STATE_TABLE1_reg_5_0_inst : FD1 port map( D => n4241, CP => CLK_I, Q => 
                           n4462, QN => n3894);
   STATE_TABLE1_reg_6_7_inst : FD1 port map( D => n4240, CP => CLK_I, Q => 
                           n4548, QN => n_3193);
   STATE_TABLE1_reg_6_6_inst : FD1 port map( D => n4239, CP => CLK_I, Q => 
                           n4437, QN => n_3194);
   STATE_TABLE1_reg_6_5_inst : FD1 port map( D => n4238, CP => CLK_I, Q => 
                           n4408, QN => n_3195);
   STATE_TABLE1_reg_6_4_inst : FD1 port map( D => n4237, CP => CLK_I, Q => 
                           n4560, QN => n_3196);
   STATE_TABLE1_reg_6_3_inst : FD1 port map( D => n4236, CP => CLK_I, Q => 
                           n4575, QN => n3889);
   STATE_TABLE1_reg_6_2_inst : FD1 port map( D => n4235, CP => CLK_I, Q => 
                           n4574, QN => n3888);
   STATE_TABLE1_reg_6_1_inst : FD1 port map( D => n4234, CP => CLK_I, Q => 
                           n4559, QN => n_3197);
   STATE_TABLE1_reg_6_0_inst : FD1 port map( D => n4233, CP => CLK_I, Q => 
                           n4573, QN => n3886);
   STATE_TABLE1_reg_7_7_inst : FD1 port map( D => n4232, CP => CLK_I, Q => 
                           n4546, QN => n_3198);
   STATE_TABLE1_reg_7_6_inst : FD1 port map( D => n4231, CP => CLK_I, Q => 
                           n4430, QN => n_3199);
   STATE_TABLE1_reg_7_5_inst : FD1 port map( D => n4230, CP => CLK_I, Q => 
                           n4528, QN => n_3200);
   STATE_TABLE1_reg_7_4_inst : FD1 port map( D => n4229, CP => CLK_I, Q => 
                           n4583, QN => n3882);
   STATE_TABLE1_reg_7_3_inst : FD1 port map( D => n4228, CP => CLK_I, Q => 
                           n4451, QN => n_3201);
   STATE_TABLE1_reg_7_2_inst : FD1 port map( D => n4227, CP => CLK_I, Q => 
                           n4582, QN => n3880);
   STATE_TABLE1_reg_7_1_inst : FD1 port map( D => n4226, CP => CLK_I, Q => 
                           n4581, QN => n3879);
   STATE_TABLE1_reg_7_0_inst : FD1 port map( D => n4225, CP => CLK_I, Q => 
                           n4429, QN => n_3202);
   STATE_TABLE1_reg_8_7_inst : FD1 port map( D => n4224, CP => CLK_I, Q => 
                           n4438, QN => n_3203);
   STATE_TABLE1_reg_8_6_inst : FD1 port map( D => n4223, CP => CLK_I, Q => 
                           n4524, QN => n_3204);
   STATE_TABLE1_reg_8_5_inst : FD1 port map( D => n4222, CP => CLK_I, Q => 
                           n4409, QN => n_3205);
   STATE_TABLE1_reg_8_4_inst : FD1 port map( D => n4221, CP => CLK_I, Q => 
                           n4594, QN => n3874);
   STATE_TABLE1_reg_8_3_inst : FD1 port map( D => n4220, CP => CLK_I, Q => 
                           n4593, QN => n3873);
   STATE_TABLE1_reg_8_2_inst : FD1 port map( D => n4219, CP => CLK_I, Q => 
                           n4592, QN => n3872);
   STATE_TABLE1_reg_8_1_inst : FD1 port map( D => n4218, CP => CLK_I, Q => 
                           n4591, QN => n3871);
   STATE_TABLE1_reg_8_0_inst : FD1 port map( D => n4217, CP => CLK_I, Q => 
                           n4590, QN => n3870);
   STATE_TABLE1_reg_9_7_inst : FD1 port map( D => n4216, CP => CLK_I, Q => 
                           n4410, QN => n_3206);
   STATE_TABLE1_reg_9_6_inst : FD1 port map( D => n4215, CP => CLK_I, Q => 
                           n4421, QN => n_3207);
   STATE_TABLE1_reg_9_5_inst : FD1 port map( D => n4214, CP => CLK_I, Q => 
                           n4597, QN => n3867);
   STATE_TABLE1_reg_9_4_inst : FD1 port map( D => n4213, CP => CLK_I, Q => 
                           n4445, QN => n_3208);
   STATE_TABLE1_reg_9_3_inst : FD1 port map( D => n4212, CP => CLK_I, Q => 
                           n4444, QN => n_3209);
   STATE_TABLE1_reg_9_2_inst : FD1 port map( D => n4211, CP => CLK_I, Q => 
                           n4383, QN => n_3210);
   STATE_TABLE1_reg_9_1_inst : FD1 port map( D => n4210, CP => CLK_I, Q => 
                           n4596, QN => n3863);
   STATE_TABLE1_reg_9_0_inst : FD1 port map( D => n4209, CP => CLK_I, Q => 
                           n4595, QN => n3862);
   STATE_TABLE1_reg_10_7_inst : FD1 port map( D => n4208, CP => CLK_I, Q => 
                           n4534, QN => n3861);
   STATE_TABLE1_reg_10_6_inst : FD1 port map( D => n4207, CP => CLK_I, Q => 
                           n4423, QN => n3860);
   STATE_TABLE1_reg_10_5_inst : FD1 port map( D => n4206, CP => CLK_I, Q => 
                           n4422, QN => n3859);
   STATE_TABLE1_reg_10_4_inst : FD1 port map( D => n4205, CP => CLK_I, Q => 
                           n4553, QN => n3858);
   STATE_TABLE1_reg_10_3_inst : FD1 port map( D => n4204, CP => CLK_I, Q => 
                           n4614, QN => n3857);
   STATE_TABLE1_reg_10_2_inst : FD1 port map( D => n4203, CP => CLK_I, Q => 
                           n4613, QN => n3856);
   STATE_TABLE1_reg_10_1_inst : FD1 port map( D => n4202, CP => CLK_I, Q => 
                           n4561, QN => n3855);
   STATE_TABLE1_reg_10_0_inst : FD1 port map( D => n4201, CP => CLK_I, Q => 
                           n4549, QN => n3854);
   STATE_TABLE1_reg_11_7_inst : FD1 port map( D => n4200, CP => CLK_I, Q => 
                           n4530, QN => n_3211);
   STATE_TABLE1_reg_11_6_inst : FD1 port map( D => n4199, CP => CLK_I, Q => 
                           n4417, QN => n_3212);
   STATE_TABLE1_reg_11_5_inst : FD1 port map( D => n4198, CP => CLK_I, Q => 
                           n4529, QN => n_3213);
   STATE_TABLE1_reg_11_4_inst : FD1 port map( D => n4197, CP => CLK_I, Q => 
                           n4469, QN => n3850);
   STATE_TABLE1_reg_11_3_inst : FD1 port map( D => n4196, CP => CLK_I, Q => 
                           n4441, QN => n_3214);
   STATE_TABLE1_reg_11_2_inst : FD1 port map( D => n4195, CP => CLK_I, Q => 
                           n4468, QN => n3848);
   STATE_TABLE1_reg_11_1_inst : FD1 port map( D => n4194, CP => CLK_I, Q => 
                           n4467, QN => n3847);
   STATE_TABLE1_reg_11_0_inst : FD1 port map( D => n4193, CP => CLK_I, Q => 
                           n4432, QN => n_3215);
   STATE_TABLE1_reg_12_7_inst : FD1 port map( D => n4192, CP => CLK_I, Q => 
                           n4446, QN => n3845);
   STATE_TABLE1_reg_12_6_inst : FD1 port map( D => n4191, CP => CLK_I, Q => 
                           n4535, QN => n3844);
   STATE_TABLE1_reg_12_5_inst : FD1 port map( D => n4190, CP => CLK_I, Q => 
                           n_3216, QN => n3843);
   STATE_TABLE1_reg_12_4_inst : FD1 port map( D => n4189, CP => CLK_I, Q => 
                           n4618, QN => n3842);
   STATE_TABLE1_reg_12_3_inst : FD1 port map( D => n4188, CP => CLK_I, Q => 
                           n4617, QN => n3841);
   STATE_TABLE1_reg_12_2_inst : FD1 port map( D => n4187, CP => CLK_I, Q => 
                           n4616, QN => n3840);
   STATE_TABLE1_reg_12_1_inst : FD1 port map( D => n4186, CP => CLK_I, Q => 
                           n4615, QN => n3839);
   STATE_TABLE1_reg_12_0_inst : FD1 port map( D => n4185, CP => CLK_I, Q => 
                           n4554, QN => n3838);
   STATE_TABLE1_reg_13_7_inst : FD1 port map( D => n4184, CP => CLK_I, Q => 
                           n4531, QN => n_3217);
   STATE_TABLE1_reg_13_6_inst : FD1 port map( D => n4183, CP => CLK_I, Q => 
                           n4382, QN => n_3218);
   STATE_TABLE1_reg_13_5_inst : FD1 port map( D => n4182, CP => CLK_I, Q => 
                           n4470, QN => n3835);
   STATE_TABLE1_reg_13_4_inst : FD1 port map( D => n4181, CP => CLK_I, Q => 
                           n4557, QN => n_3219);
   STATE_TABLE1_reg_13_3_inst : FD1 port map( D => n4180, CP => CLK_I, Q => 
                           n4388, QN => n_3220);
   STATE_TABLE1_reg_13_2_inst : FD1 port map( D => n4179, CP => CLK_I, Q => 
                           n4435, QN => n_3221);
   STATE_TABLE1_reg_13_1_inst : FD1 port map( D => n4178, CP => CLK_I, Q => 
                           n4434, QN => n_3222);
   STATE_TABLE1_reg_13_0_inst : FD1 port map( D => n4177, CP => CLK_I, Q => 
                           n4433, QN => n_3223);
   STATE_TABLE1_reg_14_7_inst : FD1 port map( D => n4176, CP => CLK_I, Q => 
                           n4589, QN => n3829);
   STATE_TABLE1_reg_14_6_inst : FD1 port map( D => n4175, CP => CLK_I, Q => 
                           n4598, QN => n3828);
   STATE_TABLE1_reg_14_5_inst : FD1 port map( D => n4174, CP => CLK_I, Q => 
                           n4541, QN => n3827);
   STATE_TABLE1_reg_14_4_inst : FD1 port map( D => n4173, CP => CLK_I, Q => 
                           n4558, QN => n_3224);
   STATE_TABLE1_reg_14_3_inst : FD1 port map( D => n4172, CP => CLK_I, Q => 
                           n4588, QN => n3825);
   STATE_TABLE1_reg_14_2_inst : FD1 port map( D => n4171, CP => CLK_I, Q => 
                           n4587, QN => n3824);
   STATE_TABLE1_reg_14_1_inst : FD1 port map( D => n4170, CP => CLK_I, Q => 
                           n4586, QN => n3823);
   STATE_TABLE1_reg_14_0_inst : FD1 port map( D => n4169, CP => CLK_I, Q => 
                           n4547, QN => n_3225);
   STATE_TABLE1_reg_15_7_inst : FD1 port map( D => n4168, CP => CLK_I, Q => 
                           n4550, QN => n3821);
   STATE_TABLE1_reg_15_6_inst : FD1 port map( D => n4167, CP => CLK_I, Q => 
                           n4424, QN => n3820);
   STATE_TABLE1_reg_15_5_inst : FD1 port map( D => n4166, CP => CLK_I, Q => 
                           n4525, QN => n3819);
   v_RAM_IN0_reg_24_inst : FD1 port map( D => n4165, CP => CLK_I, Q => n_3226, 
                           QN => n4503);
   t_STATE_RAM0_reg_0_24_inst : FD1 port map( D => n4164, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_24_port, QN => n_3227);
   t_STATE_RAM0_reg_1_24_inst : FD1 port map( D => n4163, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_24_port, QN => n_3228);
   t_STATE_RAM0_reg_2_24_inst : FD1 port map( D => n4162, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_24_port, QN => n_3229);
   t_STATE_RAM0_reg_3_24_inst : FD1 port map( D => n4161, CP => CLK_I, Q => 
                           n_3230, QN => n4665);
   v_RAM_OUT0_reg_24_inst : FD1 port map( D => n4160, CP => CLK_I, Q => 
                           v_RAM_OUT0_24_port, QN => n4374);
   STATE_TABLE1_reg_15_4_inst : FD1 port map( D => n4159, CP => CLK_I, Q => 
                           n4621, QN => n3818);
   v_RAM_IN0_reg_31_inst : FD1 port map( D => n4158, CP => CLK_I, Q => n_3231, 
                           QN => n4502);
   t_STATE_RAM0_reg_0_31_inst : FD1 port map( D => n4157, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_31_port, QN => n_3232);
   t_STATE_RAM0_reg_1_31_inst : FD1 port map( D => n4156, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_31_port, QN => n_3233);
   t_STATE_RAM0_reg_2_31_inst : FD1 port map( D => n4155, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_31_port, QN => n_3234);
   t_STATE_RAM0_reg_3_31_inst : FD1 port map( D => n4154, CP => CLK_I, Q => 
                           n_3235, QN => n4664);
   v_RAM_OUT0_reg_31_inst : FD1 port map( D => n4153, CP => CLK_I, Q => 
                           v_RAM_OUT0_31_port, QN => n4579);
   v_RAM_IN0_reg_23_inst : FD1 port map( D => n4152, CP => CLK_I, Q => n_3236, 
                           QN => n4501);
   t_STATE_RAM0_reg_0_23_inst : FD1 port map( D => n4151, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_23_port, QN => n_3237);
   t_STATE_RAM0_reg_1_23_inst : FD1 port map( D => n4150, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_23_port, QN => n_3238);
   t_STATE_RAM0_reg_2_23_inst : FD1 port map( D => n4149, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_23_port, QN => n_3239);
   t_STATE_RAM0_reg_3_23_inst : FD1 port map( D => n4148, CP => CLK_I, Q => 
                           n_3240, QN => n4663);
   v_RAM_OUT0_reg_23_inst : FD1 port map( D => n4147, CP => CLK_I, Q => 
                           v_RAM_OUT0_23_port, QN => n4564);
   v_RAM_IN0_reg_15_inst : FD1 port map( D => n4146, CP => CLK_I, Q => n_3241, 
                           QN => n4500);
   t_STATE_RAM0_reg_0_15_inst : FD1 port map( D => n4145, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_15_port, QN => n_3242);
   t_STATE_RAM0_reg_1_15_inst : FD1 port map( D => n4144, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_15_port, QN => n_3243);
   t_STATE_RAM0_reg_2_15_inst : FD1 port map( D => n4143, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_15_port, QN => n_3244);
   t_STATE_RAM0_reg_3_15_inst : FD1 port map( D => n4142, CP => CLK_I, Q => 
                           n_3245, QN => n4662);
   v_RAM_OUT0_reg_15_inst : FD1 port map( D => n4141, CP => CLK_I, Q => 
                           v_RAM_OUT0_15_port, QN => n4415);
   v_RAM_IN0_reg_7_inst : FD1 port map( D => n4140, CP => CLK_I, Q => n_3246, 
                           QN => n4499);
   t_STATE_RAM0_reg_0_7_inst : FD1 port map( D => n4139, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_7_port, QN => n_3247);
   t_STATE_RAM0_reg_1_7_inst : FD1 port map( D => n4138, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_7_port, QN => n_3248);
   t_STATE_RAM0_reg_2_7_inst : FD1 port map( D => n4137, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_7_port, QN => n_3249);
   t_STATE_RAM0_reg_3_7_inst : FD1 port map( D => n4136, CP => CLK_I, Q => 
                           n_3250, QN => n4661);
   v_RAM_OUT0_reg_7_inst : FD1 port map( D => n4135, CP => CLK_I, Q => 
                           v_RAM_OUT0_7_port, QN => n4580);
   STATE_TABLE1_reg_15_3_inst : FD1 port map( D => n4134, CP => CLK_I, Q => 
                           n4448, QN => n3817);
   v_RAM_IN0_reg_30_inst : FD1 port map( D => n4133, CP => CLK_I, Q => n_3251, 
                           QN => n4498);
   t_STATE_RAM0_reg_0_30_inst : FD1 port map( D => n4132, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_30_port, QN => n_3252);
   t_STATE_RAM0_reg_1_30_inst : FD1 port map( D => n4131, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_30_port, QN => n_3253);
   t_STATE_RAM0_reg_2_30_inst : FD1 port map( D => n4130, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_30_port, QN => n_3254);
   t_STATE_RAM0_reg_3_30_inst : FD1 port map( D => n4129, CP => CLK_I, Q => 
                           n_3255, QN => n4660);
   v_RAM_OUT0_reg_30_inst : FD1 port map( D => n4128, CP => CLK_I, Q => 
                           v_RAM_OUT0_30_port, QN => n4532);
   v_RAM_IN0_reg_22_inst : FD1 port map( D => n4127, CP => CLK_I, Q => n_3256, 
                           QN => n4497);
   t_STATE_RAM0_reg_0_22_inst : FD1 port map( D => n4126, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_22_port, QN => n_3257);
   t_STATE_RAM0_reg_1_22_inst : FD1 port map( D => n4125, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_22_port, QN => n_3258);
   t_STATE_RAM0_reg_2_22_inst : FD1 port map( D => n4124, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_22_port, QN => n_3259);
   t_STATE_RAM0_reg_3_22_inst : FD1 port map( D => n4123, CP => CLK_I, Q => 
                           n_3260, QN => n4659);
   v_RAM_OUT0_reg_22_inst : FD1 port map( D => n4122, CP => CLK_I, Q => 
                           v_RAM_OUT0_22_port, QN => n4512);
   v_RAM_IN0_reg_14_inst : FD1 port map( D => n4121, CP => CLK_I, Q => n_3261, 
                           QN => n4496);
   t_STATE_RAM0_reg_0_14_inst : FD1 port map( D => n4120, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_14_port, QN => n_3262);
   t_STATE_RAM0_reg_1_14_inst : FD1 port map( D => n4119, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_14_port, QN => n_3263);
   t_STATE_RAM0_reg_2_14_inst : FD1 port map( D => n4118, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_14_port, QN => n_3264);
   t_STATE_RAM0_reg_3_14_inst : FD1 port map( D => n4117, CP => CLK_I, Q => 
                           n_3265, QN => n4658);
   v_RAM_OUT0_reg_14_inst : FD1 port map( D => n4116, CP => CLK_I, Q => 
                           v_RAM_OUT0_14_port, QN => n4533);
   v_RAM_IN0_reg_6_inst : FD1 port map( D => n4115, CP => CLK_I, Q => n_3266, 
                           QN => n4495);
   t_STATE_RAM0_reg_0_6_inst : FD1 port map( D => n4114, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_6_port, QN => n_3267);
   t_STATE_RAM0_reg_1_6_inst : FD1 port map( D => n4113, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_6_port, QN => n_3268);
   t_STATE_RAM0_reg_2_6_inst : FD1 port map( D => n4112, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_6_port, QN => n_3269);
   t_STATE_RAM0_reg_3_6_inst : FD1 port map( D => n4111, CP => CLK_I, Q => 
                           n_3270, QN => n4657);
   v_RAM_OUT0_reg_6_inst : FD1 port map( D => n4110, CP => CLK_I, Q => 
                           v_RAM_OUT0_6_port, QN => n4511);
   STATE_TABLE1_reg_15_2_inst : FD1 port map( D => n4109, CP => CLK_I, Q => 
                           n4620, QN => n3816);
   v_RAM_IN0_reg_21_inst : FD1 port map( D => n4108, CP => CLK_I, Q => n_3271, 
                           QN => n4494);
   t_STATE_RAM0_reg_0_21_inst : FD1 port map( D => n4107, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_21_port, QN => n_3272);
   t_STATE_RAM0_reg_1_21_inst : FD1 port map( D => n4106, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_21_port, QN => n_3273);
   t_STATE_RAM0_reg_2_21_inst : FD1 port map( D => n4105, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_21_port, QN => n_3274);
   t_STATE_RAM0_reg_3_21_inst : FD1 port map( D => n4104, CP => CLK_I, Q => 
                           n_3275, QN => n4656);
   v_RAM_OUT0_reg_21_inst : FD1 port map( D => n4103, CP => CLK_I, Q => 
                           v_RAM_OUT0_21_port, QN => n4402);
   v_RAM_IN0_reg_13_inst : FD1 port map( D => n4102, CP => CLK_I, Q => n_3276, 
                           QN => n4493);
   t_STATE_RAM0_reg_0_13_inst : FD1 port map( D => n4101, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_13_port, QN => n_3277);
   t_STATE_RAM0_reg_1_13_inst : FD1 port map( D => n4100, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_13_port, QN => n_3278);
   t_STATE_RAM0_reg_2_13_inst : FD1 port map( D => n4099, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_13_port, QN => n_3279);
   t_STATE_RAM0_reg_3_13_inst : FD1 port map( D => n4098, CP => CLK_I, Q => 
                           n_3280, QN => n4655);
   v_RAM_OUT0_reg_13_inst : FD1 port map( D => n4097, CP => CLK_I, Q => 
                           v_RAM_OUT0_13_port, QN => n4519);
   v_RAM_IN0_reg_29_inst : FD1 port map( D => n4096, CP => CLK_I, Q => n_3281, 
                           QN => n4492);
   t_STATE_RAM0_reg_0_29_inst : FD1 port map( D => n4095, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_29_port, QN => n_3282);
   t_STATE_RAM0_reg_1_29_inst : FD1 port map( D => n4094, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_29_port, QN => n_3283);
   t_STATE_RAM0_reg_2_29_inst : FD1 port map( D => n4093, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_29_port, QN => n_3284);
   t_STATE_RAM0_reg_3_29_inst : FD1 port map( D => n4092, CP => CLK_I, Q => 
                           n_3285, QN => n4654);
   v_RAM_OUT0_reg_29_inst : FD1 port map( D => n4091, CP => CLK_I, Q => 
                           v_RAM_OUT0_29_port, QN => n4379);
   v_RAM_IN0_reg_5_inst : FD1 port map( D => n4090, CP => CLK_I, Q => n_3286, 
                           QN => n4491);
   t_STATE_RAM0_reg_0_5_inst : FD1 port map( D => n4089, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_5_port, QN => n_3287);
   t_STATE_RAM0_reg_1_5_inst : FD1 port map( D => n4088, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_5_port, QN => n_3288);
   t_STATE_RAM0_reg_2_5_inst : FD1 port map( D => n4087, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_5_port, QN => n_3289);
   t_STATE_RAM0_reg_3_5_inst : FD1 port map( D => n4086, CP => CLK_I, Q => 
                           n_3290, QN => n4653);
   v_RAM_OUT0_reg_5_inst : FD1 port map( D => n4085, CP => CLK_I, Q => 
                           v_RAM_OUT0_5_port, QN => n4401);
   v_RAM_IN0_reg_2_inst : FD1 port map( D => n4084, CP => CLK_I, Q => n_3291, 
                           QN => n4490);
   t_STATE_RAM0_reg_0_2_inst : FD1 port map( D => n4083, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_2_port, QN => n_3292);
   t_STATE_RAM0_reg_1_2_inst : FD1 port map( D => n4082, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_2_port, QN => n_3293);
   t_STATE_RAM0_reg_2_2_inst : FD1 port map( D => n4081, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_2_port, QN => n_3294);
   t_STATE_RAM0_reg_3_2_inst : FD1 port map( D => n4080, CP => CLK_I, Q => 
                           n_3295, QN => n4652);
   v_RAM_OUT0_reg_2_inst : FD1 port map( D => n4079, CP => CLK_I, Q => 
                           v_RAM_OUT0_2_port, QN => n4371);
   STATE_TABLE1_reg_15_1_inst : FD1 port map( D => n4078, CP => CLK_I, Q => 
                           n4619, QN => n3815);
   v_RAM_IN0_reg_18_inst : FD1 port map( D => n4077, CP => CLK_I, Q => n_3296, 
                           QN => n4489);
   t_STATE_RAM0_reg_0_18_inst : FD1 port map( D => n4076, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_18_port, QN => n_3297);
   t_STATE_RAM0_reg_1_18_inst : FD1 port map( D => n4075, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_18_port, QN => n_3298);
   t_STATE_RAM0_reg_2_18_inst : FD1 port map( D => n4074, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_18_port, QN => n_3299);
   t_STATE_RAM0_reg_3_18_inst : FD1 port map( D => n4073, CP => CLK_I, Q => 
                           n_3300, QN => n4651);
   v_RAM_OUT0_reg_18_inst : FD1 port map( D => n4072, CP => CLK_I, Q => 
                           v_RAM_OUT0_18_port, QN => n4395);
   v_RAM_IN0_reg_9_inst : FD1 port map( D => n4071, CP => CLK_I, Q => n_3301, 
                           QN => n4488);
   t_STATE_RAM0_reg_0_9_inst : FD1 port map( D => n4070, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_9_port, QN => n_3302);
   t_STATE_RAM0_reg_1_9_inst : FD1 port map( D => n4069, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_9_port, QN => n_3303);
   t_STATE_RAM0_reg_2_9_inst : FD1 port map( D => n4068, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_9_port, QN => n_3304);
   t_STATE_RAM0_reg_3_9_inst : FD1 port map( D => n4067, CP => CLK_I, Q => 
                           n_3305, QN => n4650);
   v_RAM_OUT0_reg_9_inst : FD1 port map( D => n4066, CP => CLK_I, Q => 
                           v_RAM_OUT0_9_port, QN => n4563);
   v_RAM_IN0_reg_28_inst : FD1 port map( D => n4065, CP => CLK_I, Q => n_3306, 
                           QN => n4487);
   t_STATE_RAM0_reg_0_28_inst : FD1 port map( D => n4064, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_28_port, QN => n_3307);
   t_STATE_RAM0_reg_1_28_inst : FD1 port map( D => n4063, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_28_port, QN => n_3308);
   t_STATE_RAM0_reg_2_28_inst : FD1 port map( D => n4062, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_28_port, QN => n_3309);
   t_STATE_RAM0_reg_3_28_inst : FD1 port map( D => n4061, CP => CLK_I, Q => 
                           n_3310, QN => n4649);
   v_RAM_OUT0_reg_28_inst : FD1 port map( D => n4060, CP => CLK_I, Q => 
                           v_RAM_OUT0_28_port, QN => n4359);
   v_RAM_IN0_reg_12_inst : FD1 port map( D => n4059, CP => CLK_I, Q => n_3311, 
                           QN => n4486);
   t_STATE_RAM0_reg_0_12_inst : FD1 port map( D => n4058, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_12_port, QN => n_3312);
   t_STATE_RAM0_reg_1_12_inst : FD1 port map( D => n4057, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_12_port, QN => n_3313);
   t_STATE_RAM0_reg_2_12_inst : FD1 port map( D => n4056, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_12_port, QN => n_3314);
   t_STATE_RAM0_reg_3_12_inst : FD1 port map( D => n4055, CP => CLK_I, Q => 
                           n_3315, QN => n4648);
   v_RAM_OUT0_reg_12_inst : FD1 port map( D => n4054, CP => CLK_I, Q => 
                           v_RAM_OUT0_12_port, QN => n4404);
   v_RAM_IN0_reg_20_inst : FD1 port map( D => n4053, CP => CLK_I, Q => n_3316, 
                           QN => n4485);
   t_STATE_RAM0_reg_0_20_inst : FD1 port map( D => n4052, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_20_port, QN => n_3317);
   t_STATE_RAM0_reg_1_20_inst : FD1 port map( D => n4051, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_20_port, QN => n_3318);
   t_STATE_RAM0_reg_2_20_inst : FD1 port map( D => n4050, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_20_port, QN => n_3319);
   t_STATE_RAM0_reg_3_20_inst : FD1 port map( D => n4049, CP => CLK_I, Q => 
                           n_3320, QN => n4647);
   v_RAM_OUT0_reg_20_inst : FD1 port map( D => n4048, CP => CLK_I, Q => 
                           v_RAM_OUT0_20_port, QN => n4354);
   v_RAM_IN0_reg_4_inst : FD1 port map( D => n4047, CP => CLK_I, Q => n_3321, 
                           QN => n4484);
   t_STATE_RAM0_reg_0_4_inst : FD1 port map( D => n4046, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_4_port, QN => n_3322);
   t_STATE_RAM0_reg_1_4_inst : FD1 port map( D => n4045, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_4_port, QN => n_3323);
   t_STATE_RAM0_reg_2_4_inst : FD1 port map( D => n4044, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_4_port, QN => n_3324);
   t_STATE_RAM0_reg_3_4_inst : FD1 port map( D => n4043, CP => CLK_I, Q => 
                           n_3325, QN => n4646);
   v_RAM_OUT0_reg_4_inst : FD1 port map( D => n4042, CP => CLK_I, Q => 
                           v_RAM_OUT0_4_port, QN => n4357);
   v_RAM_IN0_reg_1_inst : FD1 port map( D => n4041, CP => CLK_I, Q => n_3326, 
                           QN => n4483);
   t_STATE_RAM0_reg_0_1_inst : FD1 port map( D => n4040, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_1_port, QN => n_3327);
   t_STATE_RAM0_reg_1_1_inst : FD1 port map( D => n4039, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_1_port, QN => n_3328);
   t_STATE_RAM0_reg_2_1_inst : FD1 port map( D => n4038, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_1_port, QN => n_3329);
   t_STATE_RAM0_reg_3_1_inst : FD1 port map( D => n4037, CP => CLK_I, Q => 
                           n_3330, QN => n4645);
   v_RAM_OUT0_reg_1_inst : FD1 port map( D => n4036, CP => CLK_I, Q => 
                           v_RAM_OUT0_1_port, QN => n4508);
   STATE_TABLE1_reg_15_0_inst : FD1 port map( D => n4035, CP => CLK_I, Q => 
                           n4447, QN => n3814);
   v_RAM_IN0_reg_25_inst : FD1 port map( D => n4034, CP => CLK_I, Q => n_3331, 
                           QN => n4482);
   t_STATE_RAM0_reg_0_25_inst : FD1 port map( D => n4033, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_25_port, QN => n_3332);
   t_STATE_RAM0_reg_1_25_inst : FD1 port map( D => n4032, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_25_port, QN => n_3333);
   t_STATE_RAM0_reg_2_25_inst : FD1 port map( D => n4031, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_25_port, QN => n_3334);
   t_STATE_RAM0_reg_3_25_inst : FD1 port map( D => n4030, CP => CLK_I, Q => 
                           n_3335, QN => n4644);
   v_RAM_OUT0_reg_25_inst : FD1 port map( D => n4029, CP => CLK_I, Q => 
                           v_RAM_OUT0_25_port, QN => n4510);
   v_RAM_IN0_reg_17_inst : FD1 port map( D => n4028, CP => CLK_I, Q => n_3336, 
                           QN => n4481);
   t_STATE_RAM0_reg_0_17_inst : FD1 port map( D => n4027, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_17_port, QN => n_3337);
   t_STATE_RAM0_reg_1_17_inst : FD1 port map( D => n4026, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_17_port, QN => n_3338);
   t_STATE_RAM0_reg_2_17_inst : FD1 port map( D => n4025, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_17_port, QN => n_3339);
   t_STATE_RAM0_reg_3_17_inst : FD1 port map( D => n4024, CP => CLK_I, Q => 
                           n_3340, QN => n4643);
   v_RAM_OUT0_reg_17_inst : FD1 port map( D => n4023, CP => CLK_I, Q => 
                           v_RAM_OUT0_17_port, QN => n4509);
   v_RAM_IN0_reg_26_inst : FD1 port map( D => n4022, CP => CLK_I, Q => n_3341, 
                           QN => n4480);
   t_STATE_RAM0_reg_0_26_inst : FD1 port map( D => n4021, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_26_port, QN => n_3342);
   t_STATE_RAM0_reg_1_26_inst : FD1 port map( D => n4020, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_26_port, QN => n_3343);
   t_STATE_RAM0_reg_2_26_inst : FD1 port map( D => n4019, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_26_port, QN => n_3344);
   t_STATE_RAM0_reg_3_26_inst : FD1 port map( D => n4018, CP => CLK_I, Q => 
                           n_3345, QN => n4642);
   v_RAM_OUT0_reg_26_inst : FD1 port map( D => n4017, CP => CLK_I, Q => 
                           v_RAM_OUT0_26_port, QN => n4397);
   v_RAM_IN0_reg_10_inst : FD1 port map( D => n4016, CP => CLK_I, Q => n_3346, 
                           QN => n4479);
   t_STATE_RAM0_reg_0_10_inst : FD1 port map( D => n4015, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_10_port, QN => n_3347);
   t_STATE_RAM0_reg_1_10_inst : FD1 port map( D => n4014, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_10_port, QN => n_3348);
   t_STATE_RAM0_reg_2_10_inst : FD1 port map( D => n4013, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_10_port, QN => n_3349);
   t_STATE_RAM0_reg_3_10_inst : FD1 port map( D => n4012, CP => CLK_I, Q => 
                           n_3350, QN => n4641);
   v_RAM_OUT0_reg_10_inst : FD1 port map( D => n4011, CP => CLK_I, Q => 
                           v_RAM_OUT0_10_port, QN => n4378);
   v_RAM_IN0_reg_27_inst : FD1 port map( D => n4010, CP => CLK_I, Q => n_3351, 
                           QN => n4478);
   t_STATE_RAM0_reg_0_27_inst : FD1 port map( D => n4009, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_27_port, QN => n_3352);
   t_STATE_RAM0_reg_1_27_inst : FD1 port map( D => n4008, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_27_port, QN => n_3353);
   t_STATE_RAM0_reg_2_27_inst : FD1 port map( D => n4007, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_27_port, QN => n_3354);
   t_STATE_RAM0_reg_3_27_inst : FD1 port map( D => n4006, CP => CLK_I, Q => 
                           n_3355, QN => n4640);
   v_RAM_OUT0_reg_27_inst : FD1 port map( D => n4005, CP => CLK_I, Q => 
                           v_RAM_OUT0_27_port, QN => n4416);
   v_RAM_IN0_reg_19_inst : FD1 port map( D => n4004, CP => CLK_I, Q => n_3356, 
                           QN => n4477);
   t_STATE_RAM0_reg_0_19_inst : FD1 port map( D => n4003, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_19_port, QN => n_3357);
   t_STATE_RAM0_reg_1_19_inst : FD1 port map( D => n4002, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_19_port, QN => n_3358);
   t_STATE_RAM0_reg_2_19_inst : FD1 port map( D => n4001, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_19_port, QN => n_3359);
   t_STATE_RAM0_reg_3_19_inst : FD1 port map( D => n4000, CP => CLK_I, Q => 
                           n_3360, QN => n4639);
   v_RAM_OUT0_reg_19_inst : FD1 port map( D => n3999, CP => CLK_I, Q => 
                           v_RAM_OUT0_19_port, QN => n4399);
   v_RAM_IN0_reg_11_inst : FD1 port map( D => n3998, CP => CLK_I, Q => n_3361, 
                           QN => n4476);
   t_STATE_RAM0_reg_0_11_inst : FD1 port map( D => n3997, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_11_port, QN => n_3362);
   t_STATE_RAM0_reg_1_11_inst : FD1 port map( D => n3996, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_11_port, QN => n_3363);
   t_STATE_RAM0_reg_2_11_inst : FD1 port map( D => n3995, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_11_port, QN => n_3364);
   t_STATE_RAM0_reg_3_11_inst : FD1 port map( D => n3994, CP => CLK_I, Q => 
                           n_3365, QN => n4638);
   v_RAM_OUT0_reg_11_inst : FD1 port map( D => n3993, CP => CLK_I, Q => 
                           v_RAM_OUT0_11_port, QN => n4405);
   v_RAM_IN0_reg_3_inst : FD1 port map( D => n3992, CP => CLK_I, Q => n_3366, 
                           QN => n4475);
   t_STATE_RAM0_reg_0_3_inst : FD1 port map( D => n3991, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_3_port, QN => n_3367);
   t_STATE_RAM0_reg_1_3_inst : FD1 port map( D => n3990, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_3_port, QN => n_3368);
   t_STATE_RAM0_reg_2_3_inst : FD1 port map( D => n3989, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_3_port, QN => n_3369);
   t_STATE_RAM0_reg_3_3_inst : FD1 port map( D => n3988, CP => CLK_I, Q => 
                           n_3370, QN => n4637);
   v_RAM_OUT0_reg_3_inst : FD1 port map( D => n3987, CP => CLK_I, Q => 
                           v_RAM_OUT0_3_port, QN => n4398);
   v_RAM_IN0_reg_8_inst : FD1 port map( D => n3986, CP => CLK_I, Q => n_3371, 
                           QN => n4474);
   t_STATE_RAM0_reg_0_8_inst : FD1 port map( D => n3985, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_8_port, QN => n_3372);
   t_STATE_RAM0_reg_1_8_inst : FD1 port map( D => n3984, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_8_port, QN => n_3373);
   t_STATE_RAM0_reg_2_8_inst : FD1 port map( D => n3983, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_8_port, QN => n_3374);
   t_STATE_RAM0_reg_3_8_inst : FD1 port map( D => n3982, CP => CLK_I, Q => 
                           n_3375, QN => n4636);
   v_RAM_OUT0_reg_8_inst : FD1 port map( D => n3981, CP => CLK_I, Q => n_3376, 
                           QN => n4552);
   v_RAM_IN0_reg_16_inst : FD1 port map( D => n3980, CP => CLK_I, Q => n_3377, 
                           QN => n4473);
   t_STATE_RAM0_reg_0_16_inst : FD1 port map( D => n3979, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_16_port, QN => n_3378);
   t_STATE_RAM0_reg_1_16_inst : FD1 port map( D => n3978, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_16_port, QN => n_3379);
   t_STATE_RAM0_reg_2_16_inst : FD1 port map( D => n3977, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_16_port, QN => n_3380);
   t_STATE_RAM0_reg_3_16_inst : FD1 port map( D => n3976, CP => CLK_I, Q => 
                           n_3381, QN => n4635);
   v_RAM_OUT0_reg_16_inst : FD1 port map( D => n3975, CP => CLK_I, Q => 
                           v_RAM_OUT0_16_port, QN => n4373);
   v_RAM_IN0_reg_0_inst : FD1 port map( D => n3974, CP => CLK_I, Q => n_3382, 
                           QN => n4472);
   t_STATE_RAM0_reg_0_0_inst : FD1 port map( D => n3973, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_0_port, QN => n_3383);
   t_STATE_RAM0_reg_1_0_inst : FD1 port map( D => n3972, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_0_port, QN => n_3384);
   t_STATE_RAM0_reg_2_0_inst : FD1 port map( D => n3971, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_0_port, QN => n_3385);
   t_STATE_RAM0_reg_3_0_inst : FD1 port map( D => n3970, CP => CLK_I, Q => 
                           n_3386, QN => n4634);
   v_RAM_OUT0_reg_0_inst : FD1 port map( D => n3969, CP => CLK_I, Q => 
                           v_RAM_OUT0_0_port, QN => n4372);
   DATA_O_reg_7_inst : FD1 port map( D => n3968, CP => CLK_I, Q => 
                           DATA_O_7_port, QN => n_3387);
   DATA_O_reg_6_inst : FD1 port map( D => n3967, CP => CLK_I, Q => 
                           DATA_O_6_port, QN => n_3388);
   DATA_O_reg_5_inst : FD1 port map( D => n3966, CP => CLK_I, Q => 
                           DATA_O_5_port, QN => n_3389);
   DATA_O_reg_4_inst : FD1 port map( D => n3965, CP => CLK_I, Q => 
                           DATA_O_4_port, QN => n_3390);
   DATA_O_reg_3_inst : FD1 port map( D => n3964, CP => CLK_I, Q => 
                           DATA_O_3_port, QN => n_3391);
   DATA_O_reg_2_inst : FD1 port map( D => n3963, CP => CLK_I, Q => 
                           DATA_O_2_port, QN => n_3392);
   DATA_O_reg_1_inst : FD1 port map( D => n3962, CP => CLK_I, Q => 
                           DATA_O_1_port, QN => n_3393);
   DATA_O_reg_0_inst : FD1 port map( D => n3961, CP => CLK_I, Q => 
                           DATA_O_0_port, QN => n_3394);
   VALID_O_reg : FD1 port map( D => n3960, CP => CLK_I, Q => VALID_O, QN => 
                           n3813);
   U1248 : AN3 port map( A => n4540, B => n4380, C => n4414, Z => n1301);
   U1249 : OR3 port map( A => n5021, B => n5023, C => n1353, Z => n1349);
   U1595 : AN3 port map( A => n1461, B => n1462, C => n1463, Z => n1460);
   U1603 : OR3 port map( A => n4958, B => n4410, C => n4852, Z => n1483);
   U1607 : OR3 port map( A => n4571, B => n4421, C => n4851, Z => n1489);
   U1611 : OR3 port map( A => n4392, B => n4597, C => n4851, Z => n1494);
   U1615 : OR3 port map( A => n4963, B => n4445, C => n4851, Z => n1500);
   U1619 : OR3 port map( A => n4570, B => n4444, C => n4851, Z => n1504);
   U1623 : OR3 port map( A => n4569, B => n4383, C => n4851, Z => n1509);
   U1627 : OR3 port map( A => n4904, B => n4596, C => n4851, Z => n1514);
   U1631 : OR3 port map( A => n4391, B => n4595, C => n4851, Z => n1519);
   U1637 : OR3 port map( A => n4568, B => n4438, C => n4851, Z => n1527);
   U1641 : OR3 port map( A => n4918, B => n4524, C => n4851, Z => n1533);
   U1645 : OR3 port map( A => n4922, B => n4409, C => n4851, Z => n1537);
   U1649 : OR3 port map( A => n4461, B => n4594, C => n4851, Z => n1541);
   U1653 : OR3 port map( A => n4460, B => n4593, C => n4851, Z => n1547);
   U1657 : OR3 port map( A => n4459, B => n4592, C => n4851, Z => n1553);
   U1661 : OR3 port map( A => n4954, B => n4591, C => n4851, Z => n1559);
   U1665 : OR3 port map( A => n4968, B => n4590, C => n4851, Z => n1564);
   U1671 : OR3 port map( A => n4928, B => n4546, C => n4846, Z => n1571);
   U1675 : OR3 port map( A => n4567, B => n4430, C => n4845, Z => n1577);
   U1679 : OR3 port map( A => n4937, B => n4528, C => n4845, Z => n1582);
   U1683 : OR3 port map( A => n4390, B => n4583, C => n4845, Z => n1586);
   U1687 : OR3 port map( A => n4566, B => n4451, C => n4845, Z => n1592);
   U1691 : OR3 port map( A => n4389, B => n4582, C => n4845, Z => n1597);
   U1695 : OR3 port map( A => n4375, B => n4581, C => n4845, Z => n1603);
   U1699 : OR3 port map( A => n4565, B => n4429, C => n4845, Z => n1608);
   U1705 : OR3 port map( A => n4458, B => n4548, C => n4845, Z => n1614);
   U1709 : OR3 port map( A => n4577, B => n4437, C => n4845, Z => n1620);
   U1713 : OR3 port map( A => n4576, B => n4408, C => n4845, Z => n1625);
   U1717 : OR3 port map( A => n4953, B => n4560, C => n4845, Z => n1630);
   U1721 : OR3 port map( A => n4457, B => n4575, C => n4845, Z => n1634);
   U1727 : OR3 port map( A => n4456, B => n4574, C => n4845, Z => n1639);
   U1735 : OR3 port map( A => n4455, B => n4559, C => n4845, Z => n1665);
   U1741 : OR3 port map( A => n4454, B => n4573, C => n4845, Z => n1669);
   U1755 : OR3 port map( A => n4958, B => n4420, C => n4846, Z => n1700);
   U1759 : OR3 port map( A => n4571, B => n4384, C => n4846, Z => n1704);
   U1763 : OR3 port map( A => n4392, B => n4572, C => n4846, Z => n1707);
   U1767 : OR3 port map( A => n4963, B => n4453, C => n4846, Z => n1711);
   U1771 : OR3 port map( A => n4570, B => n4452, C => n4846, Z => n1714);
   U1775 : OR3 port map( A => n4569, B => n4436, C => n4846, Z => n1717);
   U1779 : OR3 port map( A => n4904, B => n4443, C => n4846, Z => n1720);
   U1783 : OR3 port map( A => n4391, B => n4462, C => n4846, Z => n1723);
   U1789 : OR3 port map( A => n4568, B => n4450, C => n4846, Z => n1729);
   U1794 : OR3 port map( A => n4918, B => n4539, C => n4846, Z => n1733);
   U1799 : OR3 port map( A => n4922, B => n4526, C => n4846, Z => n1736);
   U1804 : OR3 port map( A => n4461, B => n4632, C => n4846, Z => n1739);
   U1809 : OR3 port map( A => n4460, B => n4631, C => n4846, Z => n1743);
   U1814 : OR3 port map( A => n4459, B => n4630, C => n4846, Z => n1747);
   U1819 : OR3 port map( A => n4954, B => n4629, C => n4846, Z => n1751);
   U1824 : OR3 port map( A => n4968, B => n4628, C => n4846, Z => n1755);
   U1831 : OR3 port map( A => n4928, B => n4538, C => n4857, Z => n1760);
   U1836 : OR3 port map( A => n4567, B => n4427, C => n4857, Z => n1764);
   U1841 : OR3 port map( A => n4937, B => n4537, C => n4857, Z => n1767);
   U1846 : OR3 port map( A => n4390, B => n4627, C => n4857, Z => n1770);
   U1851 : OR3 port map( A => n4566, B => n4449, C => n4856, Z => n1774);
   U1856 : OR3 port map( A => n4389, B => n4626, C => n4855, Z => n1777);
   U1861 : OR3 port map( A => n4375, B => n4625, C => n4856, Z => n1781);
   U1866 : OR3 port map( A => n4565, B => n4440, C => n4855, Z => n1785);
   U1873 : OR3 port map( A => n4458, B => n4536, C => n4856, Z => n1789);
   U1878 : OR3 port map( A => n4577, B => n4426, C => n4855, Z => n1793);
   U1883 : OR3 port map( A => n4576, B => n4425, C => n4856, Z => n1796);
   U1888 : OR3 port map( A => n4953, B => n4555, C => n4857, Z => n1799);
   U1893 : OR3 port map( A => n4457, B => n4624, C => n4855, Z => n1802);
   U1898 : OR3 port map( A => n4456, B => n4623, C => n4856, Z => n1807);
   U1903 : OR3 port map( A => n4455, B => n4562, C => n4857, Z => n1811);
   U1908 : OR3 port map( A => n4454, B => n4622, C => n4855, Z => n1815);
   U1915 : OR3 port map( A => n4958, B => n4407, C => n4856, Z => n1820);
   U1919 : OR3 port map( A => n4571, B => n4419, C => n4857, Z => n1824);
   U1923 : OR3 port map( A => n4392, B => n4612, C => n4855, Z => n1827);
   U1927 : OR3 port map( A => n4963, B => n4551, C => n4856, Z => n1831);
   U1931 : OR3 port map( A => n4570, B => n4442, C => n4857, Z => n1834);
   U1935 : OR3 port map( A => n4569, B => n4418, C => n4855, Z => n1838);
   U1946 : OR3 port map( A => n4904, B => n4611, C => n4855, Z => n1860);
   U1952 : OR3 port map( A => n4391, B => n4610, C => n4856, Z => n1864);
   U1965 : OR3 port map( A => n4928, B => n4550, C => n4842, Z => n1895);
   U1970 : OR3 port map( A => n4567, B => n4424, C => n4840, Z => n1900);
   U1975 : OR3 port map( A => n4937, B => n4525, C => n4841, Z => n1903);
   U1980 : OR3 port map( A => n4390, B => n4621, C => n4840, Z => n1906);
   U1985 : OR3 port map( A => n4566, B => n4448, C => n4841, Z => n1910);
   U1990 : OR3 port map( A => n4389, B => n4620, C => n4840, Z => n1913);
   U2001 : OR3 port map( A => n4375, B => n4619, C => n4841, Z => n1936);
   U2006 : OR3 port map( A => n4565, B => n4447, C => n4840, Z => n1940);
   U2016 : AN3 port map( A => v_RAM_OUT0_25_port, B => n1954, C => n5048, Z => 
                           n1950);
   U2023 : OR3 port map( A => n4458, B => n4589, C => n4841, Z => n1969);
   U2035 : OR3 port map( A => n4953, B => n4558, C => n4840, Z => n1979);
   U2039 : OR3 port map( A => n4457, B => n4588, C => n4841, Z => n1982);
   U2043 : OR3 port map( A => n4456, B => n4587, C => n4840, Z => n1986);
   U2047 : OR3 port map( A => n4455, B => n4586, C => n4841, Z => n1990);
   U2051 : OR3 port map( A => n4454, B => n4547, C => n4840, Z => n1994);
   U2056 : OR3 port map( A => n1457, B => v_CALCULATION_CNTR_3_port, C => n5018
                           , Z => n1523);
   U2058 : OR3 port map( A => n4958, B => n4531, C => n4841, Z => n1999);
   U2092 : OR3 port map( A => n4571, B => n4382, C => n4840, Z => n2080);
   U2134 : OR3 port map( A => n4392, B => n4470, C => n4841, Z => n2150);
   U2163 : OR2 port map( A => n5145, B => n2190, Z => n2188);
   U2172 : OR3 port map( A => n4963, B => n4557, C => n4842, Z => n2202);
   U2181 : AN3 port map( A => v_RAM_OUT0_12_port, B => n4519, C => n2215, Z => 
                           n2213);
   U2193 : OR3 port map( A => n5139, B => n5123, C => n4364, Z => n2223);
   U2216 : AN3 port map( A => n2094, B => n2093, C => n5196, Z => n2250);
   U2220 : OR3 port map( A => n4570, B => n4388, C => n4840, Z => n2253);
   U2240 : OR3 port map( A => n5123, B => n5155, C => n4364, Z => n2279);
   U2264 : OR3 port map( A => n4569, B => n4435, C => n4841, Z => n2302);
   U2317 : OR3 port map( A => n4904, B => n4434, C => n4842, Z => n2341);
   U2391 : OR3 port map( A => n4391, B => n4433, C => n4840, Z => n2374);
   U2397 : OR3 port map( A => n5027, B => n2376, C => n2377, Z => n1567);
   U2416 : OR3 port map( A => n5235, B => v_RAM_OUT0_13_port, C => n1882, Z => 
                           n2387);
   U2523 : OR3 port map( A => n4568, B => n4446, C => n4841, Z => n2412);
   U2528 : OR3 port map( A => n4918, B => n4535, C => n4842, Z => n2416);
   U2537 : OR3 port map( A => n4461, B => n4618, C => n4840, Z => n2421);
   U2542 : OR3 port map( A => n4460, B => n4617, C => n4841, Z => n2425);
   U2549 : OR3 port map( A => n4459, B => n4616, C => n4842, Z => n2429);
   U2558 : OR3 port map( A => n4954, B => n4615, C => n4840, Z => n2453);
   U2565 : OR3 port map( A => n4968, B => n4554, C => n4841, Z => n2457);
   U2580 : OR3 port map( A => n4928, B => n4530, C => n4852, Z => n2485);
   U2592 : OR3 port map( A => n2507, B => n2508, C => n2509, Z => n2491);
   U2606 : AN3 port map( A => n2541, B => n2542, C => n5204, Z => n2540);
   U2618 : OR3 port map( A => n4567, B => n4417, C => n4852, Z => n2562);
   U2626 : AN3 port map( A => n2574, B => n2575, C => n2519, Z => n2573);
   U2652 : OR3 port map( A => n5074, B => n5063, C => n4728, Z => n2623);
   U2658 : OR3 port map( A => n4937, B => n4529, C => n4852, Z => n2630);
   U2698 : OR3 port map( A => n4390, B => n4469, C => n4852, Z => n2690);
   U2742 : OR3 port map( A => n4566, B => n4441, C => n4852, Z => n2737);
   U2788 : OR3 port map( A => n4389, B => n4468, C => n4852, Z => n2780);
   U2839 : OR3 port map( A => n4375, B => n4467, C => n4852, Z => n2818);
   U2899 : OR3 port map( A => n4565, B => n4432, C => n4852, Z => n2858);
   U2903 : OR3 port map( A => n5027, B => n2861, C => n2377, Z => n1674);
   U3034 : OR3 port map( A => n4458, B => n4534, C => n4852, Z => n2890);
   U3047 : OR3 port map( A => n2914, B => n2915, C => n2916, Z => n2896);
   U3061 : AN3 port map( A => n2949, B => n2950, C => n5193, Z => n2948);
   U3073 : OR3 port map( A => n4577, B => n4423, C => n4852, Z => n2968);
   U3082 : AN3 port map( A => n2981, B => n2982, C => n2927, Z => n2980);
   U3108 : OR3 port map( A => n5097, B => n5088, C => n4715, Z => n3030);
   U3114 : OR3 port map( A => n4576, B => n4422, C => n4852, Z => n3037);
   U3155 : OR3 port map( A => n4953, B => n4553, C => n4852, Z => n3098);
   U3201 : OR3 port map( A => n4457, B => n4614, C => n4852, Z => n3143);
   U3245 : OR3 port map( A => n4456, B => n4613, C => n4852, Z => n3187);
   U3303 : OR3 port map( A => n4455, B => n4561, C => n4852, Z => n3224);
   U3364 : OR3 port map( A => n4454, B => n4549, C => n4852, Z => n3263);
   U3391 : AN3 port map( A => v_RAM_OUT0_17_port, B => n1684, C => n5101, Z => 
                           n3273);
   U3495 : OR3 port map( A => n4568, B => n4431, C => n4855, Z => n3293);
   U3507 : OR3 port map( A => n3317, B => n3318, C => n3319, Z => n3299);
   U3521 : AN3 port map( A => n3352, B => n3353, C => n5206, Z => n3351);
   U3533 : OR3 port map( A => n4918, B => n4406, C => n4856, Z => n3371);
   U3541 : AN3 port map( A => n3384, B => n3385, C => n3330, Z => n3383);
   U3567 : OR3 port map( A => n5174, B => n5165, C => n4705, Z => n3433);
   U3573 : OR3 port map( A => n4922, B => n4523, C => n4855, Z => n3440);
   U3613 : OR3 port map( A => n4461, B => n4609, C => n4856, Z => n3501);
   U3658 : OR3 port map( A => n4460, B => n4608, C => n4855, Z => n3547);
   U3701 : OR3 port map( A => n4459, B => n4607, C => n4856, Z => n3591);
   U3758 : OR3 port map( A => n4954, B => n4606, C => n4855, Z => n3628);
   U3818 : OR3 port map( A => n4968, B => n4605, C => n4856, Z => n3668);
   U3847 : AN3 port map( A => v_RAM_OUT0_1_port, B => n2469, C => n5178, Z => 
                           n3681);
   U3952 : OR3 port map( A => v_CALCULATION_CNTR_3_port, B => n5027, C => n4556
                           , Z => n3699);
   U4133 : OR3 port map( A => n1457, B => v_CALCULATION_CNTR_3_port, C => n2861
                           , Z => n1342);
   U4174 : OR2 port map( A => v_CALCULATION_CNTR_7_port, B => 
                           v_CALCULATION_CNTR_6_port, Z => n3809);
   U4180 : OR3 port map( A => v_CALCULATION_CNTR_1_port, B => n5027, C => n4369
                           , Z => n3802);
   U4202 : OR3 port map( A => v_CALCULATION_CNTR_5_port, B => 
                           v_CALCULATION_CNTR_7_port, C => 
                           v_CALCULATION_CNTR_6_port, Z => n3812);
   U104 : EOI port map( A => n116, B => n117, Z => n115);
   U105 : EOI port map( A => n118, B => n119, Z => n117);
   U106 : EOI port map( A => n120, B => n121, Z => n116);
   U107 : EOI port map( A => n122, B => n123, Z => n113);
   U108 : EOI port map( A => n124, B => n125, Z => n123);
   U109 : EOI port map( A => n126, B => n127, Z => n122);
   U110 : EOI port map( A => n128, B => n129, Z => n109);
   U111 : ENI port map( A => n130, B => n131, Z => n129);
   U112 : EOI port map( A => n132, B => n133, Z => n128);
   U114 : EOI port map( A => n138, B => n139, Z => n136);
   U115 : ENI port map( A => n140, B => n141, Z => n139);
   U116 : EOI port map( A => n142, B => n143, Z => n138);
   U117 : EOI port map( A => v_KEY_COLUMN_9_port, B => v_DATA_COLUMN_9_port, Z 
                           => n135);
   U119 : AO1P port map( A => n147, B => n4370, C => n149, D => n150, Z => n146
                           );
   U120 : NR2I port map( A => n4368, B => n151, Z => n150);
   U121 : EOI port map( A => n152, B => n153, Z => n151);
   U122 : EOI port map( A => n154, B => n155, Z => n153);
   U123 : ENI port map( A => n156, B => n157, Z => n155);
   U124 : EOI port map( A => n158, B => n159, Z => n152);
   U125 : EOI port map( A => n160, B => n161, Z => n159);
   U127 : EOI port map( A => n166, B => n167, Z => n165);
   U128 : EOI port map( A => n168, B => n169, Z => n167);
   U129 : ENI port map( A => n170, B => n171, Z => n169);
   U130 : EOI port map( A => n172, B => n173, Z => n166);
   U131 : EOI port map( A => n174, B => n175, Z => n173);
   U132 : EOI port map( A => n4673, B => n4602, Z => n162);
   U133 : EOI port map( A => n177, B => n178, Z => n147);
   U134 : EOI port map( A => n179, B => n180, Z => n178);
   U135 : ENI port map( A => n181, B => n182, Z => n180);
   U136 : EOI port map( A => n183, B => n184, Z => n177);
   U137 : EOI port map( A => n185, B => n186, Z => n184);
   U143 : ENI port map( A => n199_port, B => n200_port, Z => n192_port);
   U146 : EOI port map( A => n201_port, B => n4969, Z => n197);
   U150 : EOI port map( A => n210, B => n211, Z => n209);
   U151 : ENI port map( A => n212, B => n213, Z => n211);
   U152 : EOI port map( A => n160, B => n214, Z => n210);
   U153 : EOI port map( A => n215, B => n216, Z => n208);
   U154 : ENI port map( A => n217, B => n218, Z => n216);
   U155 : EOI port map( A => n185, B => n219, Z => n215);
   U156 : EOI port map( A => n220, B => n221, Z => n206);
   U157 : EOI port map( A => n222, B => n223, Z => n221);
   U158 : EOI port map( A => n174, B => n224, Z => n220);
   U160 : EOI port map( A => n227, B => n228, Z => n226);
   U161 : ENI port map( A => n229, B => n230, Z => n228);
   U162 : EOI port map( A => n199_port, B => n231, Z => n227);
   U163 : EOI port map( A => n4672, B => v_DATA_COLUMN_7_port, Z => n225);
   U167 : EOI port map( A => n239, B => n240, Z => n238);
   U168 : EOI port map( A => n241, B => n242, Z => n239);
   U169 : EOI port map( A => n243, B => n244, Z => n242);
   U170 : EOI port map( A => n245, B => n246, Z => n237);
   U171 : EOI port map( A => n247, B => n248, Z => n245);
   U172 : EOI port map( A => n249, B => n250, Z => n248);
   U173 : EOI port map( A => n251, B => n252, Z => n235);
   U174 : EOI port map( A => n253, B => n254, Z => n251);
   U175 : EOI port map( A => n255, B => n256, Z => n254);
   U177 : EOI port map( A => n259, B => n260, Z => n258);
   U178 : EOI port map( A => n261, B => n262, Z => n260);
   U179 : EOI port map( A => n263, B => n264, Z => n259);
   U180 : EOI port map( A => v_KEY_COLUMN_6_port, B => v_DATA_COLUMN_6_port, Z 
                           => n257);
   U184 : EOI port map( A => n272, B => n273, Z => n271);
   U185 : EOI port map( A => n274, B => n275, Z => n273);
   U186 : EOI port map( A => n276, B => n277, Z => n272);
   U187 : EOI port map( A => n278, B => n279, Z => n270);
   U188 : EOI port map( A => n280, B => n281, Z => n279);
   U189 : EOI port map( A => n282, B => n283, Z => n278);
   U190 : EOI port map( A => n284, B => n285, Z => n268);
   U191 : EOI port map( A => n286, B => n287, Z => n285);
   U192 : EOI port map( A => n288, B => n289, Z => n284);
   U194 : EOI port map( A => n292, B => n293, Z => n291);
   U195 : ENI port map( A => n294, B => n295, Z => n293);
   U196 : EOI port map( A => n296, B => n297, Z => n292);
   U197 : EOI port map( A => v_KEY_COLUMN_5_port, B => v_DATA_COLUMN_5_port, Z 
                           => n290);
   U201 : EOI port map( A => n305, B => n306, Z => n304);
   U202 : EOI port map( A => n307, B => n308, Z => n306);
   U203 : EOI port map( A => n309, B => n310, Z => n305);
   U204 : EOI port map( A => n311, B => n312, Z => n303);
   U205 : EOI port map( A => n313, B => n314, Z => n312);
   U206 : EOI port map( A => n315, B => n316, Z => n311);
   U207 : EOI port map( A => n317, B => n318, Z => n301);
   U208 : EOI port map( A => n319, B => n320, Z => n318);
   U209 : EOI port map( A => n321, B => n322, Z => n317);
   U211 : EOI port map( A => n325, B => n326, Z => n324);
   U212 : EOI port map( A => n327, B => n328, Z => n326);
   U213 : EOI port map( A => n329, B => n330, Z => n325);
   U214 : EOI port map( A => n4671, B => v_DATA_COLUMN_4_port, Z => n323);
   U218 : EOI port map( A => n338, B => n339, Z => n337);
   U219 : EOI port map( A => n340, B => n341, Z => n339);
   U220 : EOI port map( A => n342, B => n343, Z => n338);
   U221 : EOI port map( A => n344, B => n345, Z => n343);
   U222 : EOI port map( A => n346, B => n347, Z => n336);
   U223 : EOI port map( A => n348, B => n349, Z => n347);
   U224 : EOI port map( A => n350, B => n351, Z => n346);
   U225 : EOI port map( A => n352, B => n353, Z => n351);
   U226 : EOI port map( A => n354, B => n355, Z => n334);
   U227 : ENI port map( A => n356, B => n357, Z => n355);
   U228 : EOI port map( A => n358, B => n359, Z => n354);
   U229 : EOI port map( A => n360, B => n361, Z => n359);
   U231 : EOI port map( A => n364, B => n365, Z => n363);
   U232 : ENI port map( A => n366, B => n367, Z => n365);
   U233 : EOI port map( A => n368, B => n369, Z => n364);
   U234 : EOI port map( A => n370, B => n371, Z => n369);
   U235 : EOI port map( A => n4670, B => v_DATA_COLUMN_3_port, Z => n362);
   U239 : EOI port map( A => n379, B => n380, Z => n378);
   U240 : EOI port map( A => n158, B => n381, Z => n379);
   U241 : EOI port map( A => n382, B => n383, Z => n377);
   U242 : EOI port map( A => n183, B => n384, Z => n382);
   U243 : EOI port map( A => n385, B => n386, Z => n375);
   U244 : EOI port map( A => n175, B => n387, Z => n385);
   U246 : EOI port map( A => n390, B => n391, Z => n389);
   U247 : EOI port map( A => n200_port, B => n392, Z => n390);
   U248 : EOI port map( A => v_KEY_COLUMN_31_port, B => v_DATA_COLUMN_31_port, 
                           Z => n388);
   U252 : EOI port map( A => n400, B => n401, Z => n399);
   U253 : EOI port map( A => n244, B => n402, Z => n400);
   U254 : EOI port map( A => n403, B => n404, Z => n402);
   U255 : EOI port map( A => n405, B => n406, Z => n398);
   U256 : EOI port map( A => n250, B => n407, Z => n405);
   U257 : EOI port map( A => n408, B => n409, Z => n407);
   U258 : EOI port map( A => n410, B => n411, Z => n396);
   U259 : EOI port map( A => n256, B => n412, Z => n410);
   U260 : EOI port map( A => n413, B => n414, Z => n412);
   U262 : EOI port map( A => n417, B => n418, Z => n416);
   U263 : EOI port map( A => n264, B => n419, Z => n417);
   U264 : EOI port map( A => n420, B => n421, Z => n419);
   U265 : EOI port map( A => n4690, B => v_DATA_COLUMN_30_port, Z => n415);
   U269 : EOI port map( A => n429, B => n430, Z => n428);
   U270 : EOI port map( A => n431, B => n432, Z => n430);
   U271 : ENI port map( A => n433, B => n434, Z => n429);
   U272 : ENI port map( A => n435, B => n436, Z => n434);
   U273 : EOI port map( A => n437, B => n438, Z => n427);
   U274 : EOI port map( A => n439, B => n440, Z => n438);
   U275 : ENI port map( A => n441, B => n442, Z => n437);
   U276 : ENI port map( A => n443, B => n444, Z => n442);
   U277 : EOI port map( A => n445, B => n446, Z => n425);
   U278 : ENI port map( A => n447, B => n448, Z => n446);
   U279 : EOI port map( A => n449, B => n450, Z => n445);
   U280 : ENI port map( A => n451, B => n452, Z => n450);
   U282 : EOI port map( A => n455, B => n456, Z => n454);
   U283 : ENI port map( A => n457, B => n458, Z => n456);
   U284 : EOI port map( A => n459, B => n460, Z => n455);
   U285 : EOI port map( A => n461, B => n462, Z => n460);
   U286 : EOI port map( A => n4669, B => v_DATA_COLUMN_2_port, Z => n453);
   U290 : EOI port map( A => n470, B => n471, Z => n469);
   U291 : EOI port map( A => n274, B => n472, Z => n471);
   U292 : EOI port map( A => n473, B => n474, Z => n274);
   U293 : EOI port map( A => n243, B => n475, Z => n470);
   U294 : EOI port map( A => n476, B => n477, Z => n468);
   U295 : EOI port map( A => n280, B => n478, Z => n477);
   U296 : EOI port map( A => n479, B => n480, Z => n280);
   U297 : EOI port map( A => n249, B => n481, Z => n476);
   U298 : EOI port map( A => n482, B => n483, Z => n466);
   U299 : EOI port map( A => n286, B => n484, Z => n483);
   U300 : EOI port map( A => n485, B => n486, Z => n286);
   U301 : EOI port map( A => n255, B => n487, Z => n482);
   U303 : EOI port map( A => n490, B => n491, Z => n489);
   U304 : EOI port map( A => n295, B => n492, Z => n491);
   U305 : EOI port map( A => n493, B => n494, Z => n295);
   U306 : EOI port map( A => n263, B => n495, Z => n490);
   U307 : EOI port map( A => v_KEY_COLUMN_29_port, B => v_DATA_COLUMN_29_port, 
                           Z => n488);
   U311 : EOI port map( A => n503, B => n504, Z => n502);
   U312 : EOI port map( A => n505, B => n506, Z => n504);
   U313 : EOI port map( A => n277, B => n310, Z => n503);
   U314 : EOI port map( A => n507, B => n508, Z => n501);
   U315 : EOI port map( A => n509, B => n510, Z => n508);
   U316 : EOI port map( A => n283, B => n316, Z => n507);
   U317 : EOI port map( A => n511, B => n512, Z => n499);
   U318 : EOI port map( A => n513, B => n514, Z => n512);
   U319 : EOI port map( A => n289, B => n322, Z => n511);
   U321 : EOI port map( A => n517, B => n518, Z => n516);
   U322 : EOI port map( A => n519, B => n520, Z => n518);
   U323 : EOI port map( A => n297, B => n330, Z => n517);
   U324 : EOI port map( A => n4689, B => v_DATA_COLUMN_28_port, Z => n515);
   U328 : EOI port map( A => n528, B => n529, Z => n527);
   U329 : EOI port map( A => n530, B => n531, Z => n529);
   U330 : EOI port map( A => n532, B => n533, Z => n528);
   U331 : EOI port map( A => n534, B => n345, Z => n533);
   U332 : EOI port map( A => n535, B => n536, Z => n526);
   U333 : EOI port map( A => n537, B => n538, Z => n536);
   U334 : EOI port map( A => n539, B => n540, Z => n535);
   U335 : EOI port map( A => n541, B => n353, Z => n540);
   U336 : EOI port map( A => n542, B => n543, Z => n524);
   U337 : EOI port map( A => n4909, B => n545, Z => n543);
   U339 : EOI port map( A => n547, B => n548, Z => n542);
   U340 : EOI port map( A => n549, B => n361, Z => n548);
   U342 : EOI port map( A => n552, B => n553, Z => n551);
   U343 : EOI port map( A => n4906, B => n555, Z => n553);
   U345 : EOI port map( A => n557, B => n558, Z => n552);
   U346 : EOI port map( A => n559, B => n371, Z => n558);
   U347 : EOI port map( A => n4688, B => v_DATA_COLUMN_27_port, Z => n550);
   U351 : EOI port map( A => n567, B => n568, Z => n566);
   U352 : EOI port map( A => n569, B => n570, Z => n568);
   U353 : EOI port map( A => n571, B => n572, Z => n567);
   U354 : EOI port map( A => n573, B => n574, Z => n565);
   U355 : EOI port map( A => n575, B => n576, Z => n574);
   U356 : EOI port map( A => n577, B => n578, Z => n573);
   U357 : EOI port map( A => n579, B => n580, Z => n563);
   U358 : ENI port map( A => n581, B => n582, Z => n580);
   U359 : EOI port map( A => n583, B => n584, Z => n579);
   U361 : EOI port map( A => n587, B => n588, Z => n586);
   U362 : EOI port map( A => n589, B => n590, Z => n588);
   U363 : EOI port map( A => n591, B => n592, Z => n587);
   U364 : EOI port map( A => n4687, B => v_DATA_COLUMN_26_port, Z => n585);
   U368 : EOI port map( A => n600, B => n601, Z => n599);
   U369 : ENI port map( A => n602, B => n603, Z => n601);
   U370 : ENI port map( A => n118, B => n435, Z => n600);
   U371 : EOI port map( A => n604, B => n605, Z => n598);
   U372 : ENI port map( A => n606, B => n607, Z => n605);
   U373 : ENI port map( A => n124, B => n443, Z => n604);
   U374 : EOI port map( A => n608, B => n609, Z => n596);
   U375 : EOI port map( A => n4925, B => n611, Z => n609);
   U377 : ENI port map( A => n130, B => n451, Z => n608);
   U379 : EOI port map( A => n615, B => n616, Z => n614);
   U380 : EOI port map( A => n4926, B => n618, Z => n616);
   U381 : EOI port map( A => n142, B => n461, Z => n615);
   U382 : EOI port map( A => n4686, B => v_DATA_COLUMN_25_port, Z => n613);
   U386 : EOI port map( A => n626, B => n627, Z => n625);
   U387 : EOI port map( A => n628, B => n629, Z => n627);
   U388 : EOI port map( A => n154, B => n630, Z => n629);
   U389 : ENI port map( A => n157, B => n631, Z => n626);
   U390 : EOI port map( A => n632, B => n633, Z => n631);
   U391 : EOI port map( A => n634, B => n635, Z => n624);
   U392 : EOI port map( A => n4910, B => n637, Z => n635);
   U393 : EOI port map( A => n179, B => n638, Z => n637);
   U395 : EOI port map( A => n182, B => n640, Z => n634);
   U396 : EOI port map( A => n641, B => n642, Z => n640);
   U397 : EOI port map( A => n643, B => n644, Z => n622);
   U398 : EOI port map( A => n645, B => n646, Z => n644);
   U399 : EOI port map( A => n168, B => n4914, Z => n646);
   U400 : ENI port map( A => n171, B => n648, Z => n643);
   U401 : EOI port map( A => n649, B => n650, Z => n648);
   U403 : EOI port map( A => n653, B => n654, Z => n652);
   U404 : EOI port map( A => n655, B => n656, Z => n654);
   U405 : EOI port map( A => n657, B => n4917, Z => n656);
   U406 : EOI port map( A => n659, B => n660, Z => n653);
   U407 : EOI port map( A => n661, B => n201_port, Z => n660);
   U408 : EOI port map( A => n4685, B => v_DATA_COLUMN_24_port, Z => n651);
   U412 : EOI port map( A => n669, B => n380, Z => n668);
   U413 : EOI port map( A => n670, B => n671, Z => n380);
   U414 : EOI port map( A => n672, B => n673, Z => n670);
   U415 : ENI port map( A => n212, B => n674, Z => n669);
   U416 : EOI port map( A => n632, B => n241, Z => n674);
   U417 : EOI port map( A => n675, B => n383, Z => n667);
   U418 : EOI port map( A => n676, B => n677, Z => n383);
   U419 : EOI port map( A => n678, B => n679, Z => n676);
   U420 : ENI port map( A => n217, B => n680, Z => n675);
   U421 : EOI port map( A => n641, B => n247, Z => n680);
   U422 : EOI port map( A => n681, B => n386, Z => n665);
   U423 : ENI port map( A => n682, B => n683, Z => n386);
   U424 : EOI port map( A => n684, B => n685, Z => n682);
   U425 : ENI port map( A => n222, B => n686, Z => n681);
   U426 : EOI port map( A => n649, B => n253, Z => n686);
   U428 : EOI port map( A => n689, B => n391, Z => n688);
   U429 : EOI port map( A => n4916, B => n691, Z => n391);
   U430 : EOI port map( A => n692, B => n4933, Z => n691);
   U431 : EOI port map( A => n229, B => n694, Z => n689);
   U432 : EOI port map( A => n661, B => n261, Z => n694);
   U433 : EOI port map( A => n4684, B => v_DATA_COLUMN_23_port, Z => n687);
   U437 : EOI port map( A => n702, B => n240, Z => n701);
   U438 : EOI port map( A => n703, B => n704, Z => n240);
   U439 : ENI port map( A => n154, B => n705, Z => n704);
   U440 : EOI port map( A => n276, B => n706, Z => n702);
   U441 : EOI port map( A => n214, B => n404, Z => n706);
   U442 : EOI port map( A => n707, B => n246, Z => n700);
   U443 : EOI port map( A => n708, B => n709, Z => n246);
   U444 : ENI port map( A => n179, B => n710, Z => n709);
   U445 : EOI port map( A => n282, B => n711, Z => n707);
   U446 : EOI port map( A => n219, B => n409, Z => n711);
   U447 : EOI port map( A => n712, B => n252, Z => n698);
   U448 : EOI port map( A => n713, B => n714, Z => n252);
   U449 : EOI port map( A => n168, B => n715, Z => n714);
   U450 : EOI port map( A => n288, B => n716, Z => n712);
   U451 : EOI port map( A => n224, B => n414, Z => n716);
   U453 : EOI port map( A => n719, B => n720, Z => n718);
   U454 : EOI port map( A => n296, B => n262, Z => n720);
   U455 : EOI port map( A => n721, B => n722, Z => n262);
   U456 : EOI port map( A => n201_port, B => n723, Z => n722);
   U457 : EOI port map( A => n231, B => n421, Z => n719);
   U458 : EOI port map( A => n4683, B => v_DATA_COLUMN_22_port, Z => n717);
   U462 : EOI port map( A => n731, B => n732, Z => n730);
   U463 : EOI port map( A => n474, B => n275, Z => n732);
   U464 : EOI port map( A => n733, B => n4934, Z => n275);
   U465 : EOI port map( A => n309, B => n735, Z => n731);
   U466 : EOI port map( A => n244, B => n475, Z => n735);
   U467 : EOI port map( A => n736, B => n737, Z => n729);
   U468 : EOI port map( A => n480, B => n281, Z => n737);
   U469 : EOI port map( A => n738, B => n4936, Z => n281);
   U470 : EOI port map( A => n315, B => n740, Z => n736);
   U471 : EOI port map( A => n250, B => n481, Z => n740);
   U472 : EOI port map( A => n741, B => n742, Z => n727);
   U473 : EOI port map( A => n486, B => n287, Z => n742);
   U474 : EOI port map( A => n743, B => n744, Z => n287);
   U475 : EOI port map( A => n321, B => n745, Z => n741);
   U476 : EOI port map( A => n256, B => n487, Z => n745);
   U478 : EOI port map( A => n748, B => n749, Z => n747);
   U479 : ENI port map( A => n294, B => n494, Z => n749);
   U480 : EOI port map( A => n750, B => n751, Z => n294);
   U481 : EOI port map( A => n329, B => n752, Z => n748);
   U482 : EOI port map( A => n264, B => n495, Z => n752);
   U483 : EOI port map( A => n4682, B => v_DATA_COLUMN_21_port, Z => n746);
   U487 : EOI port map( A => n760, B => n761, Z => n759);
   U488 : EOI port map( A => n505, B => n308, Z => n761);
   U489 : ENI port map( A => n762, B => n763, Z => n308);
   U490 : ENI port map( A => n764, B => n765, Z => n763);
   U491 : EOI port map( A => n473, B => n766, Z => n760);
   U492 : EOI port map( A => n767, B => n768, Z => n758);
   U493 : EOI port map( A => n509, B => n314, Z => n768);
   U494 : ENI port map( A => n769, B => n770, Z => n314);
   U495 : ENI port map( A => n771, B => n772, Z => n770);
   U496 : EOI port map( A => n479, B => n773, Z => n767);
   U497 : EOI port map( A => n774, B => n775, Z => n756);
   U498 : EOI port map( A => n513, B => n320, Z => n775);
   U499 : EOI port map( A => n776, B => n777, Z => n320);
   U500 : EOI port map( A => n4938, B => n779, Z => n777);
   U502 : EOI port map( A => n485, B => n781, Z => n774);
   U504 : EOI port map( A => n784, B => n785, Z => n783);
   U505 : EOI port map( A => n519, B => n328, Z => n785);
   U506 : EOI port map( A => n786, B => n787, Z => n328);
   U507 : ENI port map( A => n788, B => n789, Z => n787);
   U508 : EOI port map( A => n493, B => n790, Z => n784);
   U509 : EOI port map( A => v_KEY_COLUMN_20_port, B => v_DATA_COLUMN_20_port, 
                           Z => n782);
   U513 : EOI port map( A => n798, B => n799, Z => n797);
   U514 : EOI port map( A => n800, B => n603, Z => n799);
   U515 : ENI port map( A => n801, B => n802, Z => n603);
   U516 : ENI port map( A => n803, B => n804, Z => n802);
   U517 : EOI port map( A => n121, B => n805, Z => n798);
   U518 : EOI port map( A => n806, B => n807, Z => n796);
   U519 : EOI port map( A => n808, B => n607, Z => n807);
   U520 : ENI port map( A => n809, B => n810, Z => n607);
   U521 : ENI port map( A => n811, B => n812, Z => n810);
   U522 : EOI port map( A => n127, B => n813, Z => n806);
   U523 : EOI port map( A => n814, B => n815, Z => n794);
   U524 : EOI port map( A => n816, B => n611, Z => n815);
   U525 : EOI port map( A => n817, B => n818, Z => n611);
   U526 : ENI port map( A => n819, B => n820, Z => n818);
   U527 : EOI port map( A => n133, B => n821, Z => n814);
   U529 : EOI port map( A => n824, B => n825, Z => n823);
   U530 : EOI port map( A => n826, B => n618, Z => n825);
   U531 : EOI port map( A => n4907, B => n828, Z => n618);
   U532 : ENI port map( A => n829, B => n830, Z => n828);
   U534 : ENI port map( A => n143, B => n832, Z => n824);
   U535 : EOI port map( A => v_KEY_COLUMN_1_port, B => v_DATA_COLUMN_1_port, Z 
                           => n822);
   U539 : EOI port map( A => n840, B => n841, Z => n839);
   U540 : EOI port map( A => n340, B => n530, Z => n841);
   U541 : ENI port map( A => n842, B => n843, Z => n530);
   U542 : EOI port map( A => n844, B => n4964, Z => n843);
   U543 : ENI port map( A => n846, B => n847, Z => n340);
   U544 : EOI port map( A => n532, B => n848, Z => n840);
   U545 : EOI port map( A => n849, B => n850, Z => n848);
   U546 : EOI port map( A => n851, B => n852, Z => n838);
   U547 : EOI port map( A => n348, B => n537, Z => n852);
   U548 : ENI port map( A => n853, B => n854, Z => n537);
   U549 : EOI port map( A => n855, B => n4965, Z => n854);
   U550 : ENI port map( A => n857, B => n858, Z => n348);
   U551 : EOI port map( A => n539, B => n859, Z => n851);
   U552 : EOI port map( A => n860, B => n861, Z => n859);
   U553 : EOI port map( A => n862, B => n863, Z => n836);
   U554 : EOI port map( A => n356, B => n546, Z => n863);
   U555 : EOI port map( A => n864, B => n865, Z => n546);
   U556 : EOI port map( A => n866, B => n4966, Z => n865);
   U557 : ENI port map( A => n868, B => n869, Z => n356);
   U558 : EOI port map( A => n547, B => n870, Z => n862);
   U559 : EOI port map( A => n871, B => n872, Z => n870);
   U561 : EOI port map( A => n875, B => n876, Z => n874);
   U562 : EOI port map( A => n367, B => n555, Z => n876);
   U563 : EOI port map( A => n877, B => n878, Z => n555);
   U564 : EOI port map( A => n879, B => n4967, Z => n878);
   U565 : EOI port map( A => n881, B => n882, Z => n367);
   U566 : EOI port map( A => n557, B => n883, Z => n875);
   U567 : EOI port map( A => n884, B => n885, Z => n883);
   U568 : EOI port map( A => n4681, B => v_DATA_COLUMN_19_port, Z => n873);
   U572 : EOI port map( A => n893, B => n894, Z => n892);
   U573 : EOI port map( A => n431, B => n569, Z => n894);
   U574 : ENI port map( A => n895, B => n896, Z => n569);
   U575 : ENI port map( A => n897, B => n436, Z => n896);
   U576 : EOI port map( A => n804, B => n898, Z => n431);
   U577 : EOI port map( A => n899, B => n900, Z => n893);
   U578 : EOI port map( A => n120, B => n805, Z => n900);
   U579 : EOI port map( A => n901, B => n902, Z => n891);
   U580 : EOI port map( A => n439, B => n575, Z => n902);
   U581 : ENI port map( A => n903, B => n904, Z => n575);
   U582 : ENI port map( A => n905, B => n444, Z => n904);
   U583 : EOI port map( A => n812, B => n906, Z => n439);
   U584 : EOI port map( A => n907, B => n908, Z => n901);
   U585 : EOI port map( A => n126, B => n813, Z => n908);
   U586 : EOI port map( A => n909, B => n910, Z => n889);
   U587 : ENI port map( A => n447, B => n581, Z => n910);
   U588 : ENI port map( A => n911, B => n912, Z => n581);
   U589 : ENI port map( A => n913, B => n452, Z => n912);
   U590 : EOI port map( A => n820, B => n914, Z => n447);
   U591 : EOI port map( A => n915, B => n916, Z => n909);
   U592 : EOI port map( A => n132, B => n821, Z => n916);
   U594 : EOI port map( A => n919, B => n920, Z => n918);
   U595 : EOI port map( A => n458, B => n590, Z => n920);
   U596 : EOI port map( A => n921, B => n922, Z => n590);
   U597 : ENI port map( A => n923, B => n462, Z => n922);
   U598 : EOI port map( A => n924, B => n830, Z => n458);
   U599 : EOI port map( A => n925, B => n926, Z => n919);
   U600 : ENI port map( A => n140, B => n832, Z => n926);
   U601 : EOI port map( A => n4680, B => v_DATA_COLUMN_18_port, Z => n917);
   U605 : EOI port map( A => n934, B => n935, Z => n933);
   U606 : ENI port map( A => n602, B => n800, Z => n935);
   U607 : ENI port map( A => n119, B => n433, Z => n934);
   U608 : ENI port map( A => n571, B => n936, Z => n119);
   U609 : ENI port map( A => n803, B => n898, Z => n936);
   U610 : ENI port map( A => n937, B => n938, Z => n803);
   U611 : EOI port map( A => n939, B => n4947, Z => n938);
   U612 : EOI port map( A => n244, B => n276, Z => n939);
   U613 : EOI port map( A => n941, B => n381, Z => n937);
   U614 : EOI port map( A => n214, B => n4934, Z => n381);
   U615 : EOI port map( A => n673, B => n403, Z => n941);
   U616 : ENI port map( A => n805, B => n435, Z => n571);
   U617 : EOI port map( A => n942, B => n943, Z => n932);
   U618 : ENI port map( A => n606, B => n808, Z => n943);
   U619 : ENI port map( A => n125, B => n441, Z => n942);
   U620 : ENI port map( A => n577, B => n944, Z => n125);
   U621 : ENI port map( A => n811, B => n906, Z => n944);
   U622 : ENI port map( A => n945, B => n946, Z => n811);
   U623 : EOI port map( A => n947, B => n4949, Z => n946);
   U624 : EOI port map( A => n250, B => n282, Z => n947);
   U625 : EOI port map( A => n949, B => n384, Z => n945);
   U626 : EOI port map( A => n219, B => n4936, Z => n384);
   U627 : EOI port map( A => n679, B => n408, Z => n949);
   U628 : ENI port map( A => n813, B => n443, Z => n577);
   U629 : EOI port map( A => n950, B => n951, Z => n930);
   U630 : EOI port map( A => n816, B => n612, Z => n951);
   U631 : EOI port map( A => n131, B => n449, Z => n950);
   U632 : ENI port map( A => n583, B => n952, Z => n131);
   U633 : ENI port map( A => n819, B => n914, Z => n952);
   U634 : ENI port map( A => n953, B => n954, Z => n819);
   U635 : EOI port map( A => n955, B => n4948, Z => n954);
   U636 : EOI port map( A => n256, B => n288, Z => n955);
   U637 : EOI port map( A => n957, B => n387, Z => n953);
   U638 : EOI port map( A => n224, B => n4935, Z => n387);
   U639 : EOI port map( A => n685, B => n413, Z => n957);
   U640 : ENI port map( A => n821, B => n451, Z => n583);
   U642 : EOI port map( A => n961, B => n962, Z => n960);
   U643 : EOI port map( A => n826, B => n963, Z => n962);
   U644 : EOI port map( A => n141, B => n459, Z => n961);
   U645 : ENI port map( A => n924, B => n964, Z => n141);
   U646 : ENI port map( A => n829, B => n591, Z => n964);
   U647 : ENI port map( A => n832, B => n461, Z => n591);
   U648 : ENI port map( A => n965, B => n966, Z => n829);
   U649 : ENI port map( A => n229, B => n261, Z => n966);
   U650 : EOI port map( A => n967, B => n392, Z => n965);
   U651 : EOI port map( A => n231, B => n751, Z => n392);
   U652 : EOI port map( A => n968, B => n420, Z => n967);
   U653 : EOI port map( A => n4679, B => v_DATA_COLUMN_17_port, Z => n959);
   U655 : AO1P port map( A => n972, B => n4370, C => n973, D => n974, Z => n971
                           );
   U656 : NR2I port map( A => n4368, B => n975, Z => n974);
   U657 : EOI port map( A => n976, B => n977, Z => n975);
   U658 : EOI port map( A => n978, B => n979, Z => n977);
   U659 : ENI port map( A => n157, B => n980, Z => n976);
   U660 : EOI port map( A => n981, B => n156, Z => n980);
   U662 : EOI port map( A => n984, B => n985, Z => n983);
   U663 : EOI port map( A => n986, B => n987, Z => n985);
   U664 : ENI port map( A => n171, B => n988, Z => n984);
   U665 : EOI port map( A => n989, B => n170, Z => n988);
   U666 : EOI port map( A => n4678, B => n4601, Z => n982);
   U667 : EOI port map( A => n991, B => n992, Z => n972);
   U668 : EOI port map( A => n993, B => n994, Z => n992);
   U669 : EOI port map( A => n182, B => n995, Z => n991);
   U670 : EOI port map( A => n996, B => n181, Z => n995);
   U677 : ENI port map( A => n4920, B => n4969, Z => n1005);
   U682 : EOI port map( A => n1015, B => n1016, Z => n1014);
   U683 : EOI port map( A => n213, B => n630, Z => n1016);
   U684 : ENI port map( A => n672, B => n1017, Z => n213);
   U685 : EOI port map( A => n978, B => n4959, Z => n1017);
   U686 : EOI port map( A => n632, B => n158, Z => n978);
   U687 : EOI port map( A => n764, B => n705, Z => n672);
   U688 : EOI port map( A => n4934, B => n241, Z => n1015);
   U690 : EOI port map( A => n1020, B => n1021, Z => n1013);
   U691 : EOI port map( A => n218, B => n638, Z => n1021);
   U692 : ENI port map( A => n678, B => n1022, Z => n218);
   U693 : EOI port map( A => n4924, B => n4960, Z => n1022);
   U695 : EOI port map( A => n641, B => n4944, Z => n994);
   U696 : EOI port map( A => n771, B => n710, Z => n678);
   U697 : EOI port map( A => n4936, B => n247, Z => n1020);
   U699 : EOI port map( A => n1027, B => n1028, Z => n1011);
   U700 : EOI port map( A => n223, B => n4914, Z => n1028);
   U701 : ENI port map( A => n684, B => n1029, Z => n223);
   U702 : EOI port map( A => n986, B => n4961, Z => n1029);
   U703 : EOI port map( A => n649, B => n175, Z => n986);
   U704 : EOI port map( A => n780, B => n715, Z => n684);
   U705 : EOI port map( A => n4935, B => n253, Z => n1027);
   U708 : EOI port map( A => n1033, B => n1034, Z => n1032);
   U709 : EOI port map( A => n230, B => n4917, Z => n1034);
   U710 : ENI port map( A => n692, B => n1035, Z => n230);
   U711 : EOI port map( A => n4927, B => n4962, Z => n1035);
   U713 : ENI port map( A => n661, B => n200_port, Z => n1002);
   U714 : EOI port map( A => n788, B => n723, Z => n692);
   U715 : EOI port map( A => n751, B => n261, Z => n1033);
   U716 : EOI port map( A => v_KEY_COLUMN_15_port, B => v_DATA_COLUMN_15_port, 
                           Z => n1031);
   U720 : EOI port map( A => n1044, B => n401, Z => n1043);
   U721 : EOI port map( A => n703, B => n1045, Z => n401);
   U722 : ENI port map( A => n979, B => n764, Z => n1045);
   U723 : ENI port map( A => n277, B => n475, Z => n764);
   U724 : EOI port map( A => n733, B => n1046, Z => n703);
   U725 : EOI port map( A => n310, B => n766, Z => n733);
   U726 : ENI port map( A => n4913, B => n844, Z => n310);
   U727 : EOI port map( A => n276, B => n1048, Z => n1044);
   U728 : EOI port map( A => n673, B => n243, Z => n1048);
   U729 : EOI port map( A => n1049, B => n406, Z => n1042);
   U730 : EOI port map( A => n708, B => n1050, Z => n406);
   U731 : ENI port map( A => n993, B => n771, Z => n1050);
   U732 : ENI port map( A => n283, B => n481, Z => n771);
   U733 : EOI port map( A => n738, B => n1051, Z => n708);
   U734 : EOI port map( A => n316, B => n773, Z => n738);
   U735 : ENI port map( A => n4915, B => n855, Z => n316);
   U736 : EOI port map( A => n282, B => n1053, Z => n1049);
   U737 : EOI port map( A => n679, B => n249, Z => n1053);
   U738 : EOI port map( A => n1054, B => n411, Z => n1040);
   U739 : EOI port map( A => n713, B => n1055, Z => n411);
   U740 : EOI port map( A => n987, B => n780, Z => n1055);
   U741 : ENI port map( A => n289, B => n487, Z => n780);
   U742 : EOI port map( A => n743, B => n1056, Z => n713);
   U743 : EOI port map( A => n322, B => n781, Z => n743);
   U744 : ENI port map( A => n4914, B => n866, Z => n322);
   U745 : EOI port map( A => n288, B => n1057, Z => n1054);
   U746 : EOI port map( A => n685, B => n255, Z => n1057);
   U748 : EOI port map( A => n1060, B => n418, Z => n1059);
   U749 : EOI port map( A => n721, B => n1061, Z => n418);
   U750 : EOI port map( A => n4920, B => n788, Z => n1061);
   U751 : ENI port map( A => n297, B => n495, Z => n788);
   U752 : EOI port map( A => n750, B => n1062, Z => n721);
   U753 : EOI port map( A => n330, B => n790, Z => n750);
   U754 : ENI port map( A => n4917, B => n879, Z => n330);
   U755 : EOI port map( A => n296, B => n1063, Z => n1060);
   U756 : EOI port map( A => n968, B => n263, Z => n1063);
   U757 : EOI port map( A => n4677, B => v_DATA_COLUMN_14_port, Z => n1058);
   U761 : EOI port map( A => n1071, B => n1072, Z => n1070);
   U762 : EOI port map( A => n474, B => n472, Z => n1072);
   U763 : ENI port map( A => n1046, B => n212, Z => n472);
   U764 : EOI port map( A => n505, B => n307, Z => n1046);
   U765 : EOI port map( A => n632, B => n849, Z => n505);
   U766 : EOI port map( A => n765, B => n1073, Z => n474);
   U767 : ENI port map( A => n1074, B => n345, Z => n765);
   U768 : EOI port map( A => n630, B => n897, Z => n345);
   U769 : EOI port map( A => n850, B => n979, Z => n1074);
   U770 : EOI port map( A => n309, B => n1075, Z => n1071);
   U771 : EOI port map( A => n404, B => n277, Z => n1075);
   U772 : EOI port map( A => n4963, B => n4551, Z => n277);
   U773 : EOI port map( A => n1078, B => n1079, Z => n1069);
   U774 : EOI port map( A => n480, B => n478, Z => n1079);
   U775 : ENI port map( A => n1051, B => n217, Z => n478);
   U776 : EOI port map( A => n509, B => n313, Z => n1051);
   U777 : EOI port map( A => n641, B => n860, Z => n509);
   U778 : EOI port map( A => n772, B => n1080, Z => n480);
   U779 : ENI port map( A => n1081, B => n353, Z => n772);
   U780 : EOI port map( A => n638, B => n905, Z => n353);
   U781 : EOI port map( A => n861, B => n993, Z => n1081);
   U782 : EOI port map( A => n315, B => n1082, Z => n1078);
   U783 : EOI port map( A => n409, B => n283, Z => n1082);
   U784 : EOI port map( A => n4963, B => n4445, Z => n283);
   U785 : EOI port map( A => n1084, B => n1085, Z => n1067);
   U786 : EOI port map( A => n486, B => n484, Z => n1085);
   U787 : EOI port map( A => n1056, B => n222, Z => n484);
   U788 : EOI port map( A => n513, B => n319, Z => n1056);
   U789 : EOI port map( A => n649, B => n871, Z => n513);
   U790 : EOI port map( A => n779, B => n1086, Z => n486);
   U791 : ENI port map( A => n1087, B => n361, Z => n779);
   U792 : EOI port map( A => n1088, B => n913, Z => n361);
   U793 : EOI port map( A => n872, B => n987, Z => n1087);
   U794 : EOI port map( A => n321, B => n1089, Z => n1084);
   U795 : EOI port map( A => n414, B => n289, Z => n1089);
   U796 : EOI port map( A => n4963, B => n4453, Z => n289);
   U798 : EOI port map( A => n1093, B => n1094, Z => n1092);
   U799 : EOI port map( A => n494, B => n492, Z => n1094);
   U800 : ENI port map( A => n1062, B => n229, Z => n492);
   U801 : EOI port map( A => n519, B => n327, Z => n1062);
   U802 : EOI port map( A => n661, B => n884, Z => n519);
   U803 : EOI port map( A => n789, B => n1095, Z => n494);
   U804 : ENI port map( A => n1096, B => n371, Z => n789);
   U805 : EOI port map( A => n1097, B => n923, Z => n371);
   U806 : EOI port map( A => n885, B => n4920, Z => n1096);
   U807 : EOI port map( A => n329, B => n1098, Z => n1093);
   U808 : EOI port map( A => n421, B => n297, Z => n1098);
   U809 : EOI port map( A => n4963, B => n4557, Z => n297);
   U810 : EOI port map( A => n4676, B => v_DATA_COLUMN_13_port, Z => n1091);
   U814 : EOI port map( A => n1107, B => n1108, Z => n1106);
   U815 : EOI port map( A => n307, B => n506, Z => n1108);
   U816 : ENI port map( A => n762, B => n1109, Z => n506);
   U817 : ENI port map( A => n705, B => n1073, Z => n1109);
   U818 : ENI port map( A => n1110, B => n532, Z => n1073);
   U819 : EOI port map( A => n632, B => n899, Z => n532);
   U820 : EOI port map( A => n154, B => n342, Z => n1110);
   U821 : EOI port map( A => n4929, B => n4959, Z => n154);
   U822 : ENI port map( A => n309, B => n473, Z => n705);
   U823 : EOI port map( A => n4671, B => n3938, Z => n473);
   U824 : EOI port map( A => n4953, B => n4555, Z => n309);
   U825 : ENI port map( A => n1114, B => n1115, Z => n762);
   U826 : ENI port map( A => n847, B => n1116, Z => n1115);
   U827 : EOI port map( A => n4947, B => n120, Z => n847);
   U829 : EOI port map( A => n1117, B => n1118, Z => n1114);
   U830 : EOI port map( A => n633, B => n846, Z => n1118);
   U831 : ENI port map( A => n214, B => n435, Z => n846);
   U832 : EOI port map( A => n4954, B => n3935, Z => n435);
   U833 : ENI port map( A => n160, B => n4964, Z => n307);
   U835 : ENI port map( A => n4675, B => n4442, Z => n344);
   U836 : EOI port map( A => n475, B => n766, Z => n1107);
   U837 : EOI port map( A => n158, B => n534, Z => n766);
   U838 : EOI port map( A => n4689, B => n3914, Z => n475);
   U839 : EOI port map( A => n1121, B => n1122, Z => n1105);
   U840 : EOI port map( A => n313, B => n510, Z => n1122);
   U841 : ENI port map( A => n769, B => n1123, Z => n510);
   U842 : ENI port map( A => n710, B => n1080, Z => n1123);
   U843 : ENI port map( A => n1124, B => n539, Z => n1080);
   U844 : EOI port map( A => n641, B => n907, Z => n539);
   U845 : EOI port map( A => n179, B => n350, Z => n1124);
   U846 : EOI port map( A => n4930, B => n4960, Z => n179);
   U847 : ENI port map( A => n315, B => n479, Z => n710);
   U848 : EOI port map( A => n4671, B => n3874, Z => n479);
   U849 : EOI port map( A => n4953, B => n4553, Z => n315);
   U850 : ENI port map( A => n1127, B => n1128, Z => n769);
   U851 : ENI port map( A => n858, B => n1129, Z => n1128);
   U852 : EOI port map( A => n4949, B => n126, Z => n858);
   U854 : EOI port map( A => n1130, B => n1131, Z => n1127);
   U855 : EOI port map( A => n642, B => n857, Z => n1131);
   U856 : ENI port map( A => n219, B => n443, Z => n857);
   U857 : EOI port map( A => n4954, B => n3871, Z => n443);
   U858 : ENI port map( A => n185, B => n4965, Z => n313);
   U860 : ENI port map( A => n4675, B => n4444, Z => n352);
   U861 : EOI port map( A => n481, B => n773, Z => n1121);
   U862 : EOI port map( A => n183, B => n541, Z => n773);
   U863 : EOI port map( A => n4689, B => n3850, Z => n481);
   U864 : EOI port map( A => n1133, B => n1134, Z => n1103);
   U865 : EOI port map( A => n319, B => n514, Z => n1134);
   U866 : EOI port map( A => n776, B => n1135, Z => n514);
   U867 : ENI port map( A => n715, B => n1086, Z => n1135);
   U868 : ENI port map( A => n1136, B => n547, Z => n1086);
   U869 : EOI port map( A => n649, B => n915, Z => n547);
   U870 : EOI port map( A => n168, B => n358, Z => n1136);
   U871 : EOI port map( A => n4931, B => n4961, Z => n168);
   U872 : ENI port map( A => n321, B => n485, Z => n715);
   U873 : EOI port map( A => n4671, B => n3906, Z => n485);
   U874 : EOI port map( A => n4953, B => n4560, Z => n321);
   U875 : ENI port map( A => n1139, B => n1140, Z => n776);
   U876 : ENI port map( A => n869, B => n1141, Z => n1140);
   U877 : EOI port map( A => n4948, B => n132, Z => n869);
   U879 : EOI port map( A => n1142, B => n1143, Z => n1139);
   U880 : EOI port map( A => n650, B => n868, Z => n1143);
   U881 : ENI port map( A => n224, B => n451, Z => n868);
   U882 : EOI port map( A => n4954, B => n3903, Z => n451);
   U883 : ENI port map( A => n174, B => n4966, Z => n319);
   U885 : ENI port map( A => n4675, B => n4452, Z => n360);
   U886 : EOI port map( A => n487, B => n781, Z => n1133);
   U887 : EOI port map( A => n175, B => n549, Z => n781);
   U888 : EOI port map( A => n4689, B => n3882, Z => n487);
   U890 : EOI port map( A => n1147, B => n1148, Z => n1146);
   U891 : EOI port map( A => n327, B => n520, Z => n1148);
   U892 : EOI port map( A => n786, B => n1149, Z => n520);
   U893 : ENI port map( A => n723, B => n1095, Z => n1149);
   U894 : ENI port map( A => n1150, B => n557, Z => n1095);
   U895 : EOI port map( A => n661, B => n925, Z => n557);
   U896 : EOI port map( A => n201_port, B => n368, Z => n1150);
   U897 : EOI port map( A => n4933, B => n4962, Z => n201_port);
   U899 : ENI port map( A => n329, B => n493, Z => n723);
   U900 : EOI port map( A => n4671, B => n3842, Z => n493);
   U901 : EOI port map( A => n4953, B => n4558, Z => n329);
   U902 : ENI port map( A => n1152, B => n1153, Z => n786);
   U903 : EOI port map( A => n882, B => n1154, Z => n1153);
   U904 : EOI port map( A => n261, B => n140, Z => n882);
   U905 : EOI port map( A => n881, B => n1155, Z => n1152);
   U906 : EOI port map( A => n657, B => n1156, Z => n1155);
   U907 : ENI port map( A => n4921, B => n461, Z => n881);
   U908 : EOI port map( A => v_KEY_COLUMN_1_port, B => n3839, Z => n461);
   U909 : ENI port map( A => n199_port, B => n4967, Z => n327);
   U911 : ENI port map( A => n4675, B => n4388, Z => n370);
   U912 : EOI port map( A => n495, B => n790, Z => n1147);
   U913 : EOI port map( A => n200_port, B => n559, Z => n790);
   U914 : EOI port map( A => n4689, B => n3818, Z => n495);
   U915 : EOI port map( A => v_KEY_COLUMN_12_port, B => v_DATA_COLUMN_12_port, 
                           Z => n1145);
   U919 : EOI port map( A => n1166, B => n1167, Z => n1165);
   U920 : EOI port map( A => n341, B => n531, Z => n1167);
   U921 : ENI port map( A => n1117, B => n1116, Z => n531);
   U922 : EOI port map( A => n4929, B => n805, Z => n1116);
   U923 : EOI port map( A => n4686, B => n3911, Z => n805);
   U925 : EOI port map( A => n4959, B => n433, Z => n1117);
   U926 : ENI port map( A => n842, B => n1168, Z => n341);
   U927 : EOI port map( A => n534, B => n4939, Z => n1168);
   U929 : ENI port map( A => n4688, B => n4449, Z => n849);
   U930 : EOI port map( A => n4681, B => n3921, Z => n534);
   U931 : ENI port map( A => n1171, B => n1172, Z => n842);
   U932 : EOI port map( A => n804, B => n602, Z => n1172);
   U933 : ENI port map( A => n630, B => n157, Z => n804);
   U934 : EOI port map( A => n4968, B => n3934, Z => n157);
   U935 : EOI port map( A => n633, B => n1174, Z => n1171);
   U936 : EOI port map( A => n121, B => n898, Z => n1174);
   U937 : EOI port map( A => n158, B => n161, Z => n898);
   U938 : EOI port map( A => n342, B => n1175, Z => n1166);
   U939 : EOI port map( A => n844, B => n850, Z => n1175);
   U940 : ENI port map( A => n4943, B => n572, Z => n850);
   U942 : EOI port map( A => n4670, B => n3937, Z => n844);
   U943 : EOI port map( A => n160, B => n436, Z => n342);
   U944 : ENI port map( A => n4674, B => n4418, Z => n436);
   U945 : EOI port map( A => n1178, B => n1179, Z => n1164);
   U946 : EOI port map( A => n349, B => n538, Z => n1179);
   U947 : ENI port map( A => n1130, B => n1129, Z => n538);
   U948 : EOI port map( A => n4930, B => n813, Z => n1129);
   U949 : EOI port map( A => n4686, B => n3847, Z => n813);
   U951 : EOI port map( A => n4960, B => n441, Z => n1130);
   U952 : ENI port map( A => n853, B => n1180, Z => n349);
   U953 : EOI port map( A => n541, B => n4940, Z => n1180);
   U955 : ENI port map( A => n4688, B => n4441, Z => n860);
   U956 : EOI port map( A => n4681, B => n3857, Z => n541);
   U957 : ENI port map( A => n1183, B => n1184, Z => n853);
   U958 : EOI port map( A => n812, B => n606, Z => n1184);
   U959 : EOI port map( A => n638, B => n182, Z => n812);
   U960 : EOI port map( A => v_KEY_COLUMN_0_port, B => n3870, Z => n182);
   U961 : EOI port map( A => n642, B => n1185, Z => n1183);
   U962 : EOI port map( A => n127, B => n906, Z => n1185);
   U963 : EOI port map( A => n183, B => n186, Z => n906);
   U964 : EOI port map( A => n350, B => n1186, Z => n1178);
   U965 : EOI port map( A => n855, B => n861, Z => n1186);
   U966 : ENI port map( A => n4944, B => n578, Z => n861);
   U968 : EOI port map( A => n4670, B => n3873, Z => n855);
   U969 : EOI port map( A => n185, B => n444, Z => n350);
   U970 : ENI port map( A => n4674, B => n4383, Z => n444);
   U971 : EOI port map( A => n1188, B => n1189, Z => n1162);
   U972 : EOI port map( A => n357, B => n545, Z => n1189);
   U973 : EOI port map( A => n1142, B => n1141, Z => n545);
   U974 : EOI port map( A => n4931, B => n821, Z => n1141);
   U975 : EOI port map( A => n4686, B => n3879, Z => n821);
   U977 : EOI port map( A => n4961, B => n4905, Z => n1142);
   U978 : ENI port map( A => n864, B => n1191, Z => n357);
   U979 : EOI port map( A => n549, B => n4941, Z => n1191);
   U981 : ENI port map( A => n4688, B => n4451, Z => n871);
   U982 : EOI port map( A => n4681, B => n3889, Z => n549);
   U983 : ENI port map( A => n1194, B => n1195, Z => n864);
   U984 : EOI port map( A => n820, B => n612, Z => n1195);
   U985 : ENI port map( A => n1088, B => n171, Z => n820);
   U986 : EOI port map( A => n4968, B => n3902, Z => n171);
   U987 : EOI port map( A => n650, B => n1196, Z => n1194);
   U988 : EOI port map( A => n133, B => n914, Z => n1196);
   U989 : EOI port map( A => n175, B => n172, Z => n914);
   U990 : EOI port map( A => n358, B => n1197, Z => n1188);
   U991 : EOI port map( A => n866, B => n872, Z => n1197);
   U992 : ENI port map( A => n4945, B => n584, Z => n872);
   U994 : EOI port map( A => n4670, B => n3905, Z => n866);
   U995 : EOI port map( A => n174, B => n452, Z => n358);
   U996 : ENI port map( A => n4674, B => n4436, Z => n452);
   U998 : EOI port map( A => n1202, B => n1203, Z => n1201);
   U999 : EOI port map( A => n366, B => n556, Z => n1203);
   U1000 : EOI port map( A => n1156, B => n1154, Z => n556);
   U1001 : EOI port map( A => n968, B => n832, Z => n1154);
   U1002 : EOI port map( A => n4375, B => n3815, Z => n832);
   U1003 : EOI port map( A => n4962, B => n4908, Z => n1156);
   U1004 : ENI port map( A => n877, B => n1206, Z => n366);
   U1005 : EOI port map( A => n559, B => n4942, Z => n1206);
   U1007 : ENI port map( A => n4688, B => n4448, Z => n884);
   U1008 : EOI port map( A => n4681, B => n3825, Z => n559);
   U1009 : ENI port map( A => n1209, B => n1210, Z => n877);
   U1010 : EOI port map( A => n830, B => n963, Z => n1210);
   U1011 : ENI port map( A => n1097, B => n4969, Z => n830);
   U1013 : ENI port map( A => v_KEY_COLUMN_0_port, B => n4554, Z => n659);
   U1014 : EOI port map( A => n657, B => n1212, Z => n1209);
   U1015 : EOI port map( A => n143, B => n924, Z => n1212);
   U1016 : EOI port map( A => n200_port, B => n189, Z => n924);
   U1017 : EOI port map( A => n368, B => n1213, Z => n1202);
   U1018 : EOI port map( A => n879, B => n885, Z => n1213);
   U1019 : EOI port map( A => n200_port, B => n592, Z => n885);
   U1020 : EOI port map( A => n4670, B => n3841, Z => n879);
   U1021 : EOI port map( A => n199_port, B => n462, Z => n368);
   U1022 : ENI port map( A => n4674, B => n4435, Z => n462);
   U1023 : EOI port map( A => n4675, B => v_DATA_COLUMN_11_port, Z => n1200);
   U1027 : EOI port map( A => n1222, B => n1223, Z => n1221);
   U1028 : EOI port map( A => n570, B => n801, Z => n1223);
   U1029 : EOI port map( A => n4955, B => n433, Z => n801);
   U1030 : EOI port map( A => n4904, B => n3927, Z => n433);
   U1032 : ENI port map( A => n4679, B => n4562, Z => n120);
   U1033 : ENI port map( A => n121, B => n602, Z => n570);
   U1034 : EOI port map( A => n632, B => n1227, Z => n602);
   U1035 : EOI port map( A => n160, B => n981, Z => n121);
   U1036 : EOI port map( A => n897, B => n432, Z => n1222);
   U1037 : ENI port map( A => n895, B => n1228, Z => n432);
   U1038 : ENI port map( A => n572, B => n899, Z => n1228);
   U1039 : EOI port map( A => n4687, B => n3912, Z => n899);
   U1040 : EOI port map( A => n4680, B => n3920, Z => n572);
   U1041 : EOI port map( A => n118, B => n800, Z => n895);
   U1042 : ENI port map( A => n979, B => n1229, Z => n800);
   U1043 : EOI port map( A => n158, B => n4913, Z => n1229);
   U1045 : ENI port map( A => n4684, B => n4536, Z => n158);
   U1046 : ENI port map( A => n1231, B => n1232, Z => n118);
   U1047 : EOI port map( A => n632, B => n4959, Z => n1232);
   U1049 : ENI port map( A => n4677, B => n4419, Z => n403);
   U1050 : EOI port map( A => n4928, B => n4538, Z => n632);
   U1051 : EOI port map( A => n160, B => n673, Z => n1231);
   U1052 : ENI port map( A => n4690, B => n4427, Z => n673);
   U1053 : EOI port map( A => n4669, B => n3936, Z => n897);
   U1055 : EOI port map( A => n576, B => n809, Z => n1238);
   U1056 : EOI port map( A => n4956, B => n441, Z => n809);
   U1057 : EOI port map( A => n4904, B => n3863, Z => n441);
   U1059 : ENI port map( A => n4679, B => n4561, Z => n126);
   U1060 : ENI port map( A => n127, B => n606, Z => n576);
   U1061 : EOI port map( A => n641, B => n1241, Z => n606);
   U1062 : EOI port map( A => n185, B => n996, Z => n127);
   U1063 : EOI port map( A => n905, B => n440, Z => n1237);
   U1064 : ENI port map( A => n903, B => n1242, Z => n440);
   U1065 : ENI port map( A => n578, B => n907, Z => n1242);
   U1066 : EOI port map( A => n4687, B => n3848, Z => n907);
   U1067 : EOI port map( A => n4680, B => n3856, Z => n578);
   U1068 : EOI port map( A => n124, B => n808, Z => n903);
   U1069 : ENI port map( A => n993, B => n1243, Z => n808);
   U1070 : EOI port map( A => n183, B => n4915, Z => n1243);
   U1072 : ENI port map( A => n4684, B => n4534, Z => n183);
   U1073 : ENI port map( A => n1245, B => n1246, Z => n124);
   U1074 : EOI port map( A => n641, B => n4960, Z => n1246);
   U1076 : ENI port map( A => n4677, B => n4421, Z => n408);
   U1077 : EOI port map( A => n4928, B => n4530, Z => n641);
   U1078 : EOI port map( A => n185, B => n679, Z => n1245);
   U1079 : ENI port map( A => n4690, B => n4417, Z => n679);
   U1080 : EOI port map( A => n4669, B => n3872, Z => n905);
   U1082 : EOI port map( A => n1250, B => n1251, Z => n1218);
   U1083 : ENI port map( A => n582, B => n817, Z => n1251);
   U1084 : ENI port map( A => n132, B => n4905, Z => n817);
   U1086 : ENI port map( A => v_KEY_COLUMN_9_port, B => n4443, Z => n449);
   U1087 : ENI port map( A => n4679, B => n4559, Z => n132);
   U1088 : ENI port map( A => n133, B => n612, Z => n582);
   U1089 : EOI port map( A => n649, B => n1254, Z => n612);
   U1090 : EOI port map( A => n174, B => n989, Z => n133);
   U1091 : EOI port map( A => n913, B => n448, Z => n1250);
   U1092 : ENI port map( A => n911, B => n1255, Z => n448);
   U1093 : ENI port map( A => n584, B => n915, Z => n1255);
   U1094 : EOI port map( A => n4687, B => n3880, Z => n915);
   U1095 : EOI port map( A => n4680, B => n3888, Z => n584);
   U1096 : EOI port map( A => n130, B => n816, Z => n911);
   U1097 : ENI port map( A => n987, B => n1256, Z => n816);
   U1098 : EOI port map( A => n175, B => n4914, Z => n1256);
   U1099 : ENI port map( A => n4684, B => n4548, Z => n175);
   U1100 : ENI port map( A => n1258, B => n1259, Z => n130);
   U1101 : EOI port map( A => n649, B => n4961, Z => n1259);
   U1103 : ENI port map( A => n4677, B => n4384, Z => n413);
   U1104 : EOI port map( A => n4928, B => n4546, Z => n649);
   U1105 : EOI port map( A => n174, B => n685, Z => n1258);
   U1106 : ENI port map( A => n4690, B => n4430, Z => n685);
   U1107 : EOI port map( A => n4669, B => n3904, Z => n913);
   U1109 : EOI port map( A => n1265, B => n1266, Z => n1264);
   U1110 : EOI port map( A => n589, B => n831, Z => n1266);
   U1111 : EOI port map( A => n140, B => n4908, Z => n831);
   U1113 : ENI port map( A => v_KEY_COLUMN_9_port, B => n4434, Z => n459);
   U1114 : EOI port map( A => n4679, B => n3823, Z => n140);
   U1115 : EOI port map( A => n143, B => n4926, Z => n589);
   U1117 : EOI port map( A => n661, B => n1268, Z => n963);
   U1118 : EOI port map( A => n199_port, B => n999, Z => n143);
   U1119 : EOI port map( A => n923, B => n457, Z => n1265);
   U1120 : ENI port map( A => n921, B => n1269, Z => n457);
   U1121 : ENI port map( A => n592, B => n925, Z => n1269);
   U1122 : EOI port map( A => n4687, B => n3816, Z => n925);
   U1123 : EOI port map( A => n4680, B => n3824, Z => n592);
   U1124 : EOI port map( A => n142, B => n826, Z => n921);
   U1125 : ENI port map( A => n1270, B => n1271, Z => n826);
   U1126 : EOI port map( A => n200_port, B => n4917, Z => n1271);
   U1127 : EOI port map( A => n4684, B => n3829, Z => n200_port);
   U1128 : EOI port map( A => n231, B => n261, Z => n1270);
   U1129 : ENI port map( A => n1272, B => n1273, Z => n142);
   U1130 : EOI port map( A => n661, B => n4962, Z => n1273);
   U1132 : ENI port map( A => n4677, B => n4382, Z => n420);
   U1133 : EOI port map( A => n4928, B => n4550, Z => n661);
   U1134 : EOI port map( A => n968, B => n199_port, Z => n1272);
   U1135 : ENI port map( A => n4690, B => n4424, Z => n968);
   U1136 : EOI port map( A => n4669, B => n3840, Z => n923);
   U1137 : EOI port map( A => n4674, B => v_DATA_COLUMN_10_port, Z => n1263);
   U1140 : AO1P port map( A => n1280, B => n4370, C => n1281, D => n1282, Z => 
                           n1279);
   U1141 : NR2I port map( A => n4368, B => n1283, Z => n1282);
   U1142 : EOI port map( A => n1284, B => n1285, Z => n1283);
   U1143 : EOI port map( A => n671, B => n628, Z => n1285);
   U1144 : EOI port map( A => n981, B => n161, Z => n628);
   U1145 : EOI port map( A => n4678, B => n3918, Z => n161);
   U1146 : EOI port map( A => n4673, B => n3926, Z => n981);
   U1147 : EOI port map( A => n160, B => n630, Z => n671);
   U1148 : ENI port map( A => n4672, B => n4431, Z => n630);
   U1149 : EOI port map( A => n4958, B => n4407, Z => n160);
   U1150 : EOI port map( A => n156, B => n979, Z => n1284);
   U1151 : EOI port map( A => n214, B => n241, Z => n979);
   U1152 : ENI port map( A => n4683, B => n4426, Z => n241);
   U1153 : EOI port map( A => n4918, B => n4406, Z => n214);
   U1154 : ENI port map( A => n633, B => n1227, Z => n156);
   U1155 : EOI port map( A => n4685, B => n4440, Z => n1227);
   U1156 : EOI port map( A => n1019, B => n212, Z => n633);
   U1157 : ENI port map( A => n244, B => n276, Z => n212);
   U1158 : ENI port map( A => n4682, B => n4425, Z => n276);
   U1159 : EOI port map( A => n4922, B => n4523, Z => n244);
   U1160 : ENI port map( A => n404, B => n243, Z => n1019);
   U1161 : EOI port map( A => n4676, B => n3931, Z => n243);
   U1162 : EOI port map( A => n4937, B => n4537, Z => n404);
   U1166 : EOI port map( A => n1304, B => n1305, Z => n1303);
   U1167 : EOI port map( A => n683, B => n645, Z => n1305);
   U1168 : EOI port map( A => n989, B => n172, Z => n645);
   U1169 : EOI port map( A => n4678, B => n3886, Z => n172);
   U1170 : EOI port map( A => n4673, B => n3894, Z => n989);
   U1171 : ENI port map( A => n174, B => n4914, Z => n683);
   U1173 : ENI port map( A => n4672, B => n4450, Z => n1088);
   U1174 : EOI port map( A => n4958, B => n4420, Z => n174);
   U1175 : EOI port map( A => n170, B => n987, Z => n1304);
   U1176 : EOI port map( A => n224, B => n253, Z => n987);
   U1177 : ENI port map( A => n4683, B => n4437, Z => n253);
   U1178 : EOI port map( A => n4918, B => n4539, Z => n224);
   U1179 : ENI port map( A => n650, B => n1254, Z => n170);
   U1180 : EOI port map( A => n4685, B => n4429, Z => n1254);
   U1181 : EOI port map( A => n744, B => n222, Z => n650);
   U1182 : EOI port map( A => n256, B => n4951, Z => n222);
   U1184 : ENI port map( A => n4682, B => n4408, Z => n288);
   U1185 : EOI port map( A => n4922, B => n4526, Z => n256);
   U1186 : ENI port map( A => n414, B => n255, Z => n744);
   U1187 : EOI port map( A => n4676, B => n3899, Z => n255);
   U1188 : EOI port map( A => n4937, B => n4528, Z => n414);
   U1191 : EOI port map( A => v_KEY_COLUMN_0_port, B => n4600, Z => n1302);
   U1194 : EOI port map( A => n1319, B => n1320, Z => n1280);
   U1195 : EOI port map( A => n677, B => n639, Z => n1320);
   U1196 : ENI port map( A => n996, B => n186, Z => n639);
   U1197 : ENI port map( A => n4678, B => n4549, Z => n186);
   U1198 : EOI port map( A => n4673, B => n3862, Z => n996);
   U1199 : EOI port map( A => n185, B => n638, Z => n677);
   U1200 : ENI port map( A => n4672, B => n4438, Z => n638);
   U1201 : EOI port map( A => n4958, B => n4410, Z => n185);
   U1202 : EOI port map( A => n181, B => n993, Z => n1319);
   U1203 : EOI port map( A => n219, B => n247, Z => n993);
   U1204 : ENI port map( A => n4683, B => n4423, Z => n247);
   U1205 : EOI port map( A => n4918, B => n4524, Z => n219);
   U1206 : ENI port map( A => n642, B => n1241, Z => n181);
   U1207 : EOI port map( A => n4685, B => n4432, Z => n1241);
   U1208 : EOI port map( A => n1026, B => n217, Z => n642);
   U1209 : ENI port map( A => n250, B => n282, Z => n217);
   U1210 : ENI port map( A => n4682, B => n4422, Z => n282);
   U1211 : EOI port map( A => n4922, B => n4409, Z => n250);
   U1212 : ENI port map( A => n409, B => n249, Z => n1026);
   U1213 : EOI port map( A => n4676, B => n3867, Z => n249);
   U1214 : EOI port map( A => n4937, B => n4529, Z => n409);
   U1221 : ENI port map( A => n999, B => n4957, Z => n655);
   U1223 : ENI port map( A => n4678, B => n4547, Z => n189);
   U1224 : ENI port map( A => n4673, B => n4433, Z => n999);
   U1226 : AN2I port map( A => n4787, B => n1339, Z => n198);
   U1229 : EOI port map( A => n261, B => n4921, Z => n1336);
   U1231 : ENI port map( A => v_KEY_COLUMN_6_port, B => n4535, Z => n231);
   U1235 : ENI port map( A => n657, B => n1268, Z => n1339);
   U1236 : EOI port map( A => n4685, B => n4447, Z => n1268);
   U1237 : EOI port map( A => n229, B => n751, Z => n657);
   U1238 : EOI port map( A => n421, B => n263, Z => n751);
   U1239 : EOI port map( A => n4676, B => n3835, Z => n263);
   U1240 : EOI port map( A => n4937, B => n4525, Z => n421);
   U1241 : EOI port map( A => n264, B => n296, Z => n229);
   U1242 : EOI port map( A => n199_port, B => n4917, Z => n1330);
   U1244 : ENI port map( A => n4672, B => n4446, Z => n1097);
   U1245 : EOI port map( A => n4958, B => n4531, Z => n199_port);
   U1251 : ND2I port map( A => N203, B => n4764, Z => n1356);
   U1253 : ND2I port map( A => N202, B => n4764, Z => n1357);
   U1255 : ND2I port map( A => N201, B => n4764, Z => n1358);
   U1259 : ND2I port map( A => N199, B => n4764, Z => n1361);
   U1261 : ND2I port map( A => n4667, B => n4764, Z => n1362);
   U1297 : ND2I port map( A => n1386, B => v_CNT4_0_port, Z => n1377);
   U1333 : ND2I port map( A => n1403, B => n4380, Z => n1370);
   U1335 : ND2I port map( A => n4465, B => CE_I, Z => n1404);
   U1337 : ND2I port map( A => v_CNT4_0_port, B => n1403, Z => n1366);
   U1338 : NR2I port map( A => n4999, B => v_CNT4_1_port, Z => n1403);
   U1340 : ND2I port map( A => CE_I, B => n4380, Z => n1406);
   U1556 : ND2I port map( A => n1430, B => n4471, Z => n1435);
   U1562 : NR2I port map( A => n5005, B => n5012, Z => n1436);
   U1565 : ND2I port map( A => n5010, B => n1441, Z => n1439);
   U1573 : AO1P port map( A => n3949, B => n5013, C => n1446, D => n1426, Z => 
                           n4303);
   U1574 : NR2I port map( A => n5013, B => n3949, Z => n1426);
   U1576 : ND2I port map( A => n3959, B => VALID_DATA_I, Z => n1360);
   U1578 : NR2I port map( A => n4892, B => n3950, Z => n1424);
   U1579 : ND2I port map( A => n1448, B => n1449, Z => n4294);
   U1581 : NR2I port map( A => v_CALCULATION_CNTR_3_port, B => 
                           v_CALCULATION_CNTR_2_port, Z => n1451);
   U1586 : ND2I port map( A => n1453, B => n1454, Z => n4295);
   U1590 : ND2I port map( A => n3943, B => CE_I, Z => n103);
   U1604 : ND2I port map( A => n1485, B => n4410, Z => n1482);
   U1608 : ND2I port map( A => n1491, B => n4421, Z => n1488);
   U1612 : ND2I port map( A => n1497, B => n4597, Z => n1493);
   U1616 : ND2I port map( A => n1501, B => n4445, Z => n1499);
   U1620 : ND2I port map( A => n1506, B => n4444, Z => n1503);
   U1624 : ND2I port map( A => n1511, B => n4383, Z => n1508);
   U1628 : ND2I port map( A => n1516, B => n4596, Z => n1513);
   U1632 : ND2I port map( A => n1522, B => n4595, Z => n1518);
   U1634 : ND2I port map( A => n1486, B => n4851, Z => n1481);
   U1635 : ND2I port map( A => n4853, B => n1523, Z => n1486);
   U1638 : ND2I port map( A => n1529, B => n4438, Z => n1526);
   U1642 : ND2I port map( A => n1534, B => n4524, Z => n1532);
   U1646 : ND2I port map( A => n1538, B => n4409, Z => n1536);
   U1650 : ND2I port map( A => n1544, B => n4594, Z => n1540);
   U1654 : ND2I port map( A => n1550, B => n4593, Z => n1546);
   U1658 : ND2I port map( A => n1556, B => n4592, Z => n1552);
   U1662 : ND2I port map( A => n1561, B => n4591, Z => n1558);
   U1666 : ND2I port map( A => n1566, B => n4590, Z => n1563);
   U1668 : ND2I port map( A => n4759, B => n4853, Z => n1525);
   U1669 : ND2I port map( A => n4852, B => n1567, Z => n1530);
   U1672 : ND2I port map( A => n1573, B => n4546, Z => n1570);
   U1676 : ND2I port map( A => n1579, B => n4430, Z => n1576);
   U1680 : ND2I port map( A => n1583, B => n4528, Z => n1581);
   U1684 : ND2I port map( A => n1589, B => n4583, Z => n1585);
   U1688 : ND2I port map( A => n1594, B => n4451, Z => n1591);
   U1692 : ND2I port map( A => n1600, B => n4582, Z => n1596);
   U1696 : ND2I port map( A => n1605, B => n4581, Z => n1602);
   U1700 : ND2I port map( A => n1610, B => n4429, Z => n1607);
   U1702 : ND2I port map( A => n1574, B => n4845, Z => n1569);
   U1703 : ND2I port map( A => n4847, B => n1567, Z => n1574);
   U1706 : ND2I port map( A => n1616, B => n4548, Z => n1613);
   U1710 : ND2I port map( A => n1622, B => n4437, Z => n1619);
   U1714 : ND2I port map( A => n1627, B => n4408, Z => n1624);
   U1718 : ND2I port map( A => n1631, B => n4560, Z => n1629);
   U1722 : ND2I port map( A => n1637, B => n4575, Z => n1633);
   U1725 : ND2I port map( A => n1641, B => n4574, Z => n1640);
   U1731 : ND2I port map( A => n1654, B => n1655, Z => n1653);
   U1736 : ND2I port map( A => n1667, B => n4559, Z => n1664);
   U1739 : ND2I port map( A => n1671, B => n4573, Z => n1670);
   U1742 : ND2I port map( A => n4757, B => n4847, Z => n1612);
   U1743 : ND2I port map( A => n4846, B => n1674, Z => n1617);
   U1756 : ND2I port map( A => n1701, B => n4420, Z => n1699);
   U1760 : ND2I port map( A => n1705, B => n4384, Z => n1703);
   U1764 : ND2I port map( A => n1709, B => n4572, Z => n1706);
   U1768 : ND2I port map( A => n1712, B => n4453, Z => n1710);
   U1772 : ND2I port map( A => n1715, B => n4452, Z => n1713);
   U1776 : ND2I port map( A => n1718, B => n4436, Z => n1716);
   U1780 : ND2I port map( A => n1721, B => n4443, Z => n1719);
   U1784 : ND2I port map( A => n1725, B => n4462, Z => n1722);
   U1786 : ND2I port map( A => n4755, B => n4846, Z => n1698);
   U1787 : ND2I port map( A => n4846, B => n1726, Z => n1702);
   U1790 : ND2I port map( A => n1730, B => n4450, Z => n1728);
   U1795 : ND2I port map( A => n1734, B => n4539, Z => n1732);
   U1800 : ND2I port map( A => n1737, B => n4526, Z => n1735);
   U1805 : ND2I port map( A => n1741, B => n4632, Z => n1738);
   U1810 : ND2I port map( A => n1745, B => n4631, Z => n1742);
   U1815 : ND2I port map( A => n1749, B => n4630, Z => n1746);
   U1820 : ND2I port map( A => n1753, B => n4629, Z => n1750);
   U1825 : ND2I port map( A => n1757, B => n4628, Z => n1754);
   U1828 : ND2I port map( A => n4753, B => n4846, Z => n1727);
   U1829 : ND2I port map( A => n4846, B => n1523, Z => n1731);
   U1832 : ND2I port map( A => n1761, B => n4538, Z => n1759);
   U1837 : ND2I port map( A => n1765, B => n4427, Z => n1763);
   U1842 : ND2I port map( A => n1768, B => n4537, Z => n1766);
   U1847 : ND2I port map( A => n1772, B => n4627, Z => n1769);
   U1852 : ND2I port map( A => n1775, B => n4449, Z => n1773);
   U1857 : ND2I port map( A => n1779, B => n4626, Z => n1776);
   U1862 : ND2I port map( A => n1783, B => n4625, Z => n1780);
   U1867 : ND2I port map( A => n1786, B => n4440, Z => n1784);
   U1870 : ND2I port map( A => n4751, B => n4856, Z => n1758);
   U1871 : ND2I port map( A => n4857, B => n1523, Z => n1762);
   U1874 : ND2I port map( A => n1790, B => n4536, Z => n1788);
   U1879 : ND2I port map( A => n1794, B => n4426, Z => n1792);
   U1884 : ND2I port map( A => n1797, B => n4425, Z => n1795);
   U1889 : ND2I port map( A => n1800, B => n4555, Z => n1798);
   U1894 : ND2I port map( A => n1804, B => n4624, Z => n1801);
   U1899 : ND2I port map( A => n1809, B => n4623, Z => n1806);
   U1904 : ND2I port map( A => n1812, B => n4562, Z => n1810);
   U1909 : ND2I port map( A => n1817, B => n4622, Z => n1814);
   U1912 : ND2I port map( A => n4749, B => n4857, Z => n1787);
   U1913 : ND2I port map( A => n4857, B => n1567, Z => n1791);
   U1916 : ND2I port map( A => n1821, B => n4407, Z => n1819);
   U1920 : ND2I port map( A => n1825, B => n4419, Z => n1823);
   U1924 : ND2I port map( A => n1829, B => n4612, Z => n1826);
   U1928 : ND2I port map( A => n1832, B => n4551, Z => n1830);
   U1932 : ND2I port map( A => n1835, B => n4442, Z => n1833);
   U1936 : ND2I port map( A => n1839, B => n4418, Z => n1837);
   U1941 : ND2I port map( A => n5149, B => n5196, Z => n1848);
   U1943 : AO1P port map( A => n5197, B => n1854, C => n1855, D => n1856, Z => 
                           n1852);
   U1944 : NR2I port map( A => n1857, B => n1858, Z => n1855);
   U1947 : ND2I port map( A => n1862, B => n4611, Z => n1859);
   U1950 : ND2I port map( A => n1866, B => n4610, Z => n1865);
   U1953 : ND2I port map( A => n4747, B => n4855, Z => n1818);
   U1954 : ND2I port map( A => n4857, B => n1674, Z => n1822);
   U1958 : ND2I port map( A => n1879, B => n4519, Z => n1878);
   U1966 : ND2I port map( A => n1897, B => n4550, Z => n1894);
   U1971 : ND2I port map( A => n1901, B => n4424, Z => n1899);
   U1976 : ND2I port map( A => n1904, B => n4525, Z => n1902);
   U1981 : ND2I port map( A => n1908, B => n4621, Z => n1905);
   U1986 : ND2I port map( A => n1911, B => n4448, Z => n1909);
   U1991 : ND2I port map( A => n1915, B => n4620, Z => n1912);
   U1997 : AO1P port map( A => n5075, B => n1926, C => n1927, D => n1928, Z => 
                           n1923);
   U1998 : NR2I port map( A => n4838, B => n1930, Z => n1928);
   U2002 : ND2I port map( A => n1938, B => n4619, Z => n1935);
   U2007 : ND2I port map( A => n1941, B => n4447, Z => n1939);
   U2010 : ND2I port map( A => n4745, B => n4842, Z => n1893);
   U2011 : ND2I port map( A => n4842, B => n1726, Z => n1898);
   U2014 : AO1P port map( A => n5228, B => n1949, C => n1950, D => n1951, Z => 
                           n1945);
   U2015 : AN2I port map( A => n5230, B => n1953, Z => n1951);
   U2024 : ND2I port map( A => n1971, B => n4589, Z => n1968);
   U2029 : EOI port map( A => n4683, B => n3828, Z => n261);
   U2033 : ENI port map( A => n4682, B => n4541, Z => n296);
   U2036 : ND2I port map( A => n1980, B => n4558, Z => n1978);
   U2040 : ND2I port map( A => n1984, B => n4588, Z => n1981);
   U2044 : ND2I port map( A => n1988, B => n4587, Z => n1985);
   U2048 : ND2I port map( A => n1992, B => n4586, Z => n1989);
   U2052 : ND2I port map( A => n1995, B => n4547, Z => n1993);
   U2054 : ND2I port map( A => n4743, B => n4841, Z => n1967);
   U2055 : ND2I port map( A => n4842, B => n1523, Z => n1972);
   U2060 : ND2I port map( A => n2000, B => n4531, Z => n1998);
   U2066 : NR2I port map( A => v_RAM_OUT0_12_port, B => n4552, Z => n2010);
   U2072 : NR2I port map( A => v_RAM_OUT0_12_port, B => n4519, Z => n2030);
   U2081 : NR2I port map( A => n2053, B => n2054, Z => n2042);
   U2084 : AO1P port map( A => n5143, B => n5201, C => n2062, D => n2063, Z => 
                           n2040);
   U2086 : ND2I port map( A => n2068, B => n2069, Z => n2067);
   U2088 : ND2I port map( A => n2072, B => n2073, Z => n2046);
   U2089 : AO1P port map( A => n5197, B => n5142, C => n2075, D => n4415, Z => 
                           n2039);
   U2094 : ND2I port map( A => n2081, B => n4382, Z => n2079);
   U2099 : AO1P port map( A => n4766, B => n2033, C => n2091, D => n2092, Z => 
                           n2090);
   U2100 : NR2I port map( A => n4413, B => n2093, Z => n2092);
   U2104 : AO1P port map( A => n5152, B => n4767, C => n5116, D => n2101, Z => 
                           n2098);
   U2106 : ND2I port map( A => n5151, B => n4769, Z => n2097);
   U2114 : NR2I port map( A => v_RAM_OUT0_10_port, B => n4519, Z => n2117);
   U2115 : AO1P port map( A => v_RAM_OUT0_15_port, B => n2121, C => n2122, D =>
                           n2123, Z => n2082);
   U2118 : ND2I port map( A => n2129, B => n2120, Z => n2128);
   U2119 : ND2I port map( A => n2093, B => n2068, Z => n2127);
   U2127 : ND2I port map( A => n1889, B => n2021, Z => n2142);
   U2131 : AN2I port map( A => n2146, B => n2130, Z => n2034);
   U2136 : ND2I port map( A => n2152, B => n4470, Z => n2149);
   U2139 : AO1P port map( A => v_RAM_OUT0_15_port, B => n2155, C => n2156, D =>
                           n2157, Z => n2154);
   U2140 : NR2I port map( A => n2158, B => n4740, Z => n2157);
   U2141 : AO1P port map( A => n5118, B => n4766, C => n2160, D => n2161, Z => 
                           n2158);
   U2145 : AO1P port map( A => n2165, B => n4767, C => n2166, D => n2167, Z => 
                           n2156);
   U2153 : ND2I port map( A => n2072, B => n2140, Z => n2077);
   U2154 : AO1P port map( A => n4387, B => n2175, C => n2176, D => n2177, Z => 
                           n2153);
   U2155 : AO1P port map( A => n1890, B => n4765, C => n2178, D => n2179, Z => 
                           n2177);
   U2157 : NR2I port map( A => n5145, B => n5120, Z => n2180);
   U2160 : ND2I port map( A => n2184, B => n4519, Z => n2183);
   U2165 : AO1P port map( A => n4515, B => n1884, C => n2192, D => n2193, Z => 
                           n2181);
   U2166 : NR2I port map( A => n4376, B => n2194, Z => n2193);
   U2168 : ND2I port map( A => n2197, B => n2198, Z => n2175);
   U2174 : ND2I port map( A => n2203, B => n4557, Z => n2201);
   U2176 : ND2I port map( A => n2204, B => n2205, Z => n1498);
   U2178 : ND2I port map( A => v_RAM_OUT0_15_port, B => n2209, Z => n2208);
   U2182 : ND2I port map( A => n2195, B => n5199, Z => n2211);
   U2183 : NR2I port map( A => n5117, B => n1854, Z => n2195);
   U2184 : ND2I port map( A => n2216, B => n2015, Z => n2173);
   U2186 : ND2I port map( A => n2219, B => n2220, Z => n2218);
   U2188 : NR2I port map( A => n5136, B => n2215, Z => n2165);
   U2194 : ND2I port map( A => n2094, B => n2093, Z => n2222);
   U2196 : NR2I port map( A => n5116, B => n2230, Z => n2229);
   U2201 : AO1P port map( A => n5072, B => n2236, C => n5069, D => 
                           v_RAM_OUT0_9_port, Z => n2235);
   U2207 : ND2I port map( A => n5125, B => n2112, Z => n2133);
   U2210 : ND2I port map( A => n5117, B => n4770, Z => n2231);
   U2222 : ND2I port map( A => n2254, B => n4388, Z => n2252);
   U2226 : AO1P port map( A => n2050, B => n5203, C => n2261, D => n2262, Z => 
                           n2260);
   U2228 : NR2I port map( A => n5120, B => n5136, Z => n2263);
   U2230 : NR2I port map( A => n2021, B => n5130, Z => n2050);
   U2231 : AO1P port map( A => n5241, B => n5197, C => n2267, D => n2268, Z => 
                           n2259);
   U2233 : AO1P port map( A => n5199, B => n2270, C => n2271, D => n2272, Z => 
                           n2258);
   U2236 : ND2I port map( A => n2275, B => n5125, Z => n2270);
   U2237 : AO1P port map( A => n5198, B => n2111, C => n1844, D => n2276, Z => 
                           n2257);
   U2238 : AO1P port map( A => n4515, B => n5153, C => n2277, D => n4519, Z => 
                           n2276);
   U2241 : ND2I port map( A => n4766, B => n2281, Z => n2278);
   U2244 : AO1P port map( A => n4768, B => n2194, C => n2286, D => n2287, Z => 
                           n2285);
   U2245 : NR2I port map( A => n4412, B => n2094, Z => n2287);
   U2247 : ND2I port map( A => n2275, B => n5141, Z => n2194);
   U2252 : ND2I port map( A => n2094, B => n2291, Z => n2281);
   U2256 : ND2I port map( A => n2069, B => n2214, Z => n2297);
   U2257 : NR2I port map( A => n5134, B => n5155, Z => n2296);
   U2260 : ND2I port map( A => n2072, B => n2129, Z => n2189);
   U2266 : ND2I port map( A => n2303, B => n4435, Z => n2301);
   U2269 : ND2I port map( A => n5067, B => n1845, Z => n2305);
   U2272 : ND2I port map( A => n2275, B => n2130, Z => n2312);
   U2273 : ND2I port map( A => n2164, B => n2120, Z => n2311);
   U2275 : ND2I port map( A => n2291, B => n2143, Z => n2313);
   U2277 : ND2I port map( A => n2146, B => n2120, Z => n2111);
   U2279 : ND2I port map( A => n2072, B => n2214, Z => n2264);
   U2280 : ND2I port map( A => n2164, B => n4405, Z => n2269);
   U2286 : ND2I port map( A => n4767, B => n2320, Z => n2317);
   U2287 : ND2I port map( A => n2196, B => n2143, Z => n2225);
   U2290 : ND2I port map( A => n4378, B => n4519, Z => n1857);
   U2292 : ND2I port map( A => n2214, B => n2196, Z => n2321);
   U2293 : ND2I port map( A => n2095, B => n2140, Z => n2057);
   U2297 : AO1P port map( A => n5197, B => n2214, C => n2330, D => n4415, Z => 
                           n2329);
   U2300 : ND2I port map( A => n2094, B => n5125, Z => n2135);
   U2301 : ND2I port map( A => n5196, B => n2130, Z => n2327);
   U2302 : ND2I port map( A => n5147, B => n4552, Z => n2130);
   U2304 : ND2I port map( A => n2070, B => n2116, Z => n2334);
   U2305 : NR2I port map( A => v_RAM_OUT0_13_port, B => n4404, Z => n2332);
   U2307 : AO1P port map( A => n4769, B => n2337, C => n2230, D => n2338, Z => 
                           n2336);
   U2309 : ND2I port map( A => n2072, B => n2146, Z => n2337);
   U2312 : AO1P port map( A => n4504, B => n2199, C => n2339, D => n2230, Z => 
                           n2323);
   U2313 : NR2I port map( A => n2291, B => n4365, Z => n2230);
   U2315 : NR2I port map( A => n5145, B => n2215, Z => n2018);
   U2319 : ND2I port map( A => n2342, B => n4434, Z => n2340);
   U2323 : AO1P port map( A => n5146, B => n5201, C => n2350, D => n2351, Z => 
                           n2348);
   U2325 : NR2I port map( A => n5123, B => n5148, Z => n2119);
   U2329 : ND2I port map( A => n2072, B => n1889, Z => n2023);
   U2333 : NR2I port map( A => n5144, B => n5154, Z => n2265);
   U2335 : ND2I port map( A => n2055, B => n5197, Z => n2346);
   U2337 : ND2I port map( A => n4415, B => n4563, Z => n1844);
   U2339 : ND2I port map( A => n2110, B => n5199, Z => n2354);
   U2341 : NR2I port map( A => n5240, B => n5152, Z => n2110);
   U2349 : ND2I port map( A => n2214, B => n2021, Z => n2358);
   U2350 : NR2I port map( A => n5117, B => n2190, Z => n2059);
   U2353 : ND2I port map( A => v_RAM_OUT0_15_port, B => n4563, Z => n2268);
   U2356 : AO1P port map( A => n4765, B => n2363, C => n2364, D => n2365, Z => 
                           n2362);
   U2359 : NR2I port map( A => n5144, B => n2215, Z => n2055);
   U2360 : NR2I port map( A => n5147, B => n4777, Z => n2215);
   U2361 : AO1P port map( A => n5153, B => n4768, C => n2366, D => n2191, Z => 
                           n2361);
   U2363 : ND2I port map( A => n2214, B => n2093, Z => n2367);
   U2365 : ND2I port map( A => n2072, B => n2143, Z => n2035);
   U2366 : NR2I port map( A => n5241, B => n5133, Z => n2319);
   U2370 : ND2I port map( A => n4770, B => v_RAM_OUT0_13_port, Z => n2066);
   U2372 : ND2I port map( A => n4766, B => v_RAM_OUT0_13_port, Z => n2116);
   U2375 : ND2I port map( A => n4768, B => v_RAM_OUT0_13_port, Z => n2065);
   U2377 : ND2I port map( A => n5140, B => n2164, Z => n2145);
   U2378 : ND2I port map( A => n4778, B => n2069, Z => n2164);
   U2380 : ND2I port map( A => n4769, B => v_RAM_OUT0_13_port, Z => n2109);
   U2381 : ND2I port map( A => n5197, B => n2012, Z => n2369);
   U2382 : ND2I port map( A => n2273, B => n2196, Z => n2012);
   U2385 : ND2I port map( A => n4515, B => n4519, Z => n2078);
   U2387 : NR2I port map( A => n2190, B => n5139, Z => n2251);
   U2389 : ND2I port map( A => n5140, B => n4771, Z => n2143);
   U2393 : ND2I port map( A => n2375, B => n4433, Z => n2373);
   U2395 : ND2I port map( A => n4741, B => n4842, Z => n1997);
   U2396 : ND2I port map( A => n4842, B => n1567, Z => n2001);
   U2405 : ND2I port map( A => n2068, B => n2095, Z => n2320);
   U2406 : ND2I port map( A => n4772, B => n2033, Z => n2068);
   U2408 : ND2I port map( A => v_RAM_OUT0_14_port, B => n4775, Z => n2129);
   U2410 : ND2I port map( A => n2214, B => n2095, Z => n2384);
   U2413 : ND2I port map( A => n5197, B => n2168, Z => n2388);
   U2414 : ND2I port map( A => n1889, B => n2069, Z => n2168);
   U2417 : ND2I port map( A => n2095, B => n2146, Z => n1882);
   U2418 : ND2I port map( A => n5123, B => n4776, Z => n2146);
   U2419 : ND2I port map( A => n2073, B => n2196, Z => n1884);
   U2420 : ND2I port map( A => n2021, B => n4552, Z => n2196);
   U2421 : ND2I port map( A => n4777, B => n4533, Z => n2073);
   U2424 : NR2I port map( A => n1854, B => n5133, Z => n1890);
   U2426 : ND2I port map( A => n4365, B => n4739, Z => n1881);
   U2429 : ND2I port map( A => n2291, B => n2112, Z => n2200);
   U2432 : NR2I port map( A => n5143, B => n5155, Z => n2391);
   U2434 : ND2I port map( A => n4778, B => n2162, Z => n2214);
   U2436 : ND2I port map( A => n4552, B => n2093, Z => n2216);
   U2440 : ND2I port map( A => n2401, B => n2402, Z => n2400);
   U2442 : ND2I port map( A => n4771, B => n2021, Z => n2094);
   U2444 : ND2I port map( A => n1889, B => n2120, Z => n2298);
   U2445 : ND2I port map( A => n2033, B => n4552, Z => n2120);
   U2448 : ND2I port map( A => n4519, B => n4415, Z => n2044);
   U2449 : ND2I port map( A => n2403, B => n2404, Z => n2399);
   U2453 : NR2I port map( A => n5120, B => n5133, Z => n2148);
   U2456 : ND2I port map( A => n4533, B => n4552, Z => n2291);
   U2458 : ND2I port map( A => n2095, B => n2273, Z => n2071);
   U2459 : ND2I port map( A => n5147, B => n4772, Z => n2273);
   U2461 : ND2I port map( A => v_RAM_OUT0_14_port, B => n4405, Z => n2069);
   U2462 : ND2I port map( A => v_RAM_OUT0_14_port, B => n4552, Z => n2095);
   U2465 : ND2I port map( A => v_RAM_OUT0_13_port, B => v_RAM_OUT0_15_port, Z 
                           => n2182);
   U2467 : AO1P port map( A => n4768, B => n2363, C => n2406, D => n1856, Z => 
                           n2405);
   U2468 : NR2I port map( A => n2140, B => n4378, Z => n1856);
   U2469 : ND2I port map( A => n5153, B => n4773, Z => n2140);
   U2470 : NR2I port map( A => n4737, B => n2199, Z => n2406);
   U2471 : ND2I port map( A => n2275, B => n2241, Z => n2199);
   U2472 : ND2I port map( A => n2162, B => n4552, Z => n2241);
   U2473 : ND2I port map( A => n4774, B => n4405, Z => n2275);
   U2474 : ND2I port map( A => n2015, B => n2032, Z => n2363);
   U2475 : ND2I port map( A => n5153, B => n4552, Z => n2032);
   U2476 : ND2I port map( A => n5134, B => n4771, Z => n2015);
   U2479 : ND2I port map( A => v_RAM_OUT0_13_port, B => n4415, Z => n1876);
   U2480 : ND2I port map( A => v_RAM_OUT0_10_port, B => v_RAM_OUT0_12_port, Z 
                           => n2056);
   U2482 : ND2I port map( A => n4552, B => n4405, Z => n2072);
   U2489 : ND2I port map( A => n4507, B => n4519, Z => n2210);
   U2491 : ND2I port map( A => v_RAM_OUT0_10_port, B => n4404, Z => n2102);
   U2493 : NR2I port map( A => n2033, B => n4772, Z => n2394);
   U2495 : ND2I port map( A => v_RAM_OUT0_10_port, B => n4519, Z => n2274);
   U2497 : NR2I port map( A => n1854, B => n5242, Z => n1888);
   U2498 : NR2I port map( A => n2021, B => n4773, Z => n1854);
   U2499 : ND2I port map( A => n2093, B => n2162, Z => n2021);
   U2500 : NR2I port map( A => n5153, B => n5136, Z => n2134);
   U2502 : ND2I port map( A => n4774, B => n2093, Z => n1889);
   U2504 : ND2I port map( A => v_RAM_OUT0_11_port, B => v_RAM_OUT0_14_port, Z 
                           => n2162);
   U2506 : ND2I port map( A => n4504, B => n4519, Z => n2070);
   U2508 : ND2I port map( A => v_RAM_OUT0_12_port, B => n4378, Z => n2049);
   U2509 : NR2I port map( A => n2190, B => n5242, Z => n2147);
   U2511 : ND2I port map( A => v_RAM_OUT0_11_port, B => n4773, Z => n2112);
   U2512 : NR2I port map( A => n2093, B => n4774, Z => n2190);
   U2513 : ND2I port map( A => n4533, B => n4405, Z => n2093);
   U2516 : ND2I port map( A => n4506, B => n4519, Z => n2076);
   U2519 : ND2I port map( A => n4378, B => n4404, Z => n2060);
   U2524 : ND2I port map( A => n2413, B => n4446, Z => n2411);
   U2529 : ND2I port map( A => n2417, B => n4535, Z => n2415);
   U2535 : EOI port map( A => v_KEY_COLUMN_5_port, B => n3843, Z => n264);
   U2538 : ND2I port map( A => n2423, B => n4618, Z => n2420);
   U2543 : ND2I port map( A => n2427, B => n4617, Z => n2424);
   U2547 : ND2I port map( A => n2431, B => n4616, Z => n2430);
   U2554 : ND2I port map( A => n2443, B => n2444, Z => n2442);
   U2559 : ND2I port map( A => n2455, B => n4615, Z => n2452);
   U2563 : ND2I port map( A => n2459, B => n4554, Z => n2458);
   U2567 : ND2I port map( A => n4734, B => n4840, Z => n2410);
   U2568 : ND2I port map( A => n4842, B => n1674, Z => n2414);
   U2582 : ND2I port map( A => n2486, B => n4530, Z => n2484);
   U2596 : NR2I port map( A => n4397, B => n4510, Z => n2517);
   U2605 : AO1P port map( A => n5205, B => n5076, C => n2539, D => n2540, Z => 
                           n2528);
   U2613 : ND2I port map( A => n2521, B => n2553, Z => n2501);
   U2620 : ND2I port map( A => n2563, B => n4417, Z => n2561);
   U2625 : AO1P port map( A => n2571, B => n4510, C => n2572, D => n2573, Z => 
                           n2570);
   U2628 : ND2I port map( A => n5038, B => n2581, Z => n2571);
   U2634 : ND2I port map( A => n5051, B => n4397, Z => n2592);
   U2637 : ND2I port map( A => n2597, B => n2598, Z => n2552);
   U2639 : ND2I port map( A => n2601, B => n2602, Z => n2565);
   U2641 : AO1P port map( A => n5231, B => n5074, C => n2607, D => n2608, Z => 
                           n2604);
   U2642 : NR2I port map( A => n4828, B => n2575, Z => n2608);
   U2645 : AO1P port map( A => n4833, B => n2614, C => n2615, D => n2616, Z => 
                           n2613);
   U2647 : NR2I port map( A => n5075, B => n4725, Z => n2615);
   U2653 : AO1P port map( A => n5234, B => n2625, C => n2626, D => n2627, Z => 
                           n2619);
   U2656 : ND2I port map( A => n2618, B => n1930, Z => n2625);
   U2660 : ND2I port map( A => n2631, B => n4529, Z => n2629);
   U2664 : NR2I port map( A => n2636, B => n2637, Z => n2635);
   U2673 : AO1P port map( A => n4832, B => n2550, C => v_RAM_OUT0_25_port, D =>
                           n2654, Z => n2653);
   U2674 : NR2I port map( A => n4726, B => n2609, Z => n2654);
   U2678 : NR2I port map( A => n4781, B => n5034, Z => n2659);
   U2679 : ND2I port map( A => v_RAM_OUT0_31_port, B => n2662, Z => n2634);
   U2681 : AO1P port map( A => n5231, B => n2665, C => n2666, D => n2667, Z => 
                           n2664);
   U2684 : ND2I port map( A => n2574, B => n2534, Z => n2665);
   U2694 : AO1P port map( A => n5057, B => n5231, C => n2685, D => n2686, Z => 
                           n2671);
   U2696 : NR2I port map( A => n5046, B => n5057, Z => n2556);
   U2700 : ND2I port map( A => n2692, B => n4469, Z => n2689);
   U2702 : ND2I port map( A => n2693, B => n2694, Z => n1584);
   U2711 : ND2I port map( A => n2534, B => n2708, Z => n2677);
   U2712 : NR2I port map( A => n5055, B => n5047, Z => n2683);
   U2714 : NR2I port map( A => v_RAM_OUT0_29_port, B => n4828, Z => n2703);
   U2718 : ND2I port map( A => n2657, B => n2610, Z => n2700);
   U2722 : NR2I port map( A => n2714, B => n4725, Z => n2686);
   U2727 : NR2I port map( A => n5029, B => n5058, Z => n2722);
   U2734 : AO1P port map( A => n5231, B => n2728, C => n2729, D => n2730, Z => 
                           n2727);
   U2737 : ND2I port map( A => n2534, B => n2553, Z => n2728);
   U2744 : ND2I port map( A => n2738, B => n4441, Z => n2736);
   U2749 : ND2I port map( A => n2746, B => n2747, Z => n2745);
   U2754 : ND2I port map( A => n5234, B => n2657, Z => n2750);
   U2757 : ND2I port map( A => n5075, B => n2541, Z => n2559);
   U2761 : ND2I port map( A => n2521, B => n2732, Z => n2758);
   U2763 : ND2I port map( A => n2609, B => n2708, Z => n2761);
   U2764 : NR2I port map( A => n5074, B => n5060, Z => n2760);
   U2765 : NR2I port map( A => n5060, B => n5077, Z => n2755);
   U2768 : AO1P port map( A => n4830, B => n2682, C => n2766, D => n2767, Z => 
                           n2765);
   U2769 : NR2I port map( A => n4726, B => n2610, Z => n2767);
   U2771 : ND2I port map( A => n2499, B => n2516, Z => n2682);
   U2772 : AO1P port map( A => n5032, B => n5234, C => n2769, D => n2770, Z => 
                           n2764);
   U2775 : NR2I port map( A => n5051, B => n5056, Z => n2593);
   U2777 : AO1P port map( A => n5078, B => n5232, C => n2774, D => n2775, Z => 
                           n2772);
   U2778 : NR2I port map( A => n5060, B => n2776, Z => n2775);
   U2780 : AO1P port map( A => n4827, B => n2777, C => n1962, D => n4510, Z => 
                           n2774);
   U2781 : ND2I port map( A => n2778, B => n4397, Z => n2777);
   U2783 : ND2I port map( A => n2731, B => n2610, Z => n2778);
   U2784 : ND2I port map( A => n2609, B => n1930, Z => n1933);
   U2786 : ND2I port map( A => n2782, B => n4468, Z => n2781);
   U2796 : ND2I port map( A => n2521, B => n2668, Z => n2754);
   U2802 : ND2I port map( A => n2499, B => n2598, Z => n2795);
   U2804 : ND2I port map( A => n2796, B => n2597, Z => n2585);
   U2805 : NR2I port map( A => n5054, B => n5032, Z => n2748);
   U2808 : ND2I port map( A => n2579, B => n2707, Z => n2525);
   U2810 : NR2I port map( A => n2799, B => n2800, Z => n2786);
   U2813 : ND2I port map( A => n2752, B => n2574, Z => n2649);
   U2814 : NR2I port map( A => n5063, B => n5032, Z => n2735);
   U2818 : ND2I port map( A => n2804, B => n2805, Z => n2803);
   U2826 : ND2I port map( A => n5077, B => n4374, Z => n2598);
   U2828 : ND2I port map( A => n4835, B => n2575, Z => n2807);
   U2831 : ND2I port map( A => n4724, B => n2669, Z => n2814);
   U2832 : ND2I port map( A => v_RAM_OUT0_27_port, B => n4374, Z => n2669);
   U2834 : ND2I port map( A => n2618, B => n2610, Z => n2614);
   U2835 : AN2I port map( A => n2684, B => n2793, Z => n2701);
   U2841 : ND2I port map( A => n2820, B => n4467, Z => n2817);
   U2848 : ND2I port map( A => n2499, B => n2628, Z => n2600);
   U2853 : ND2I port map( A => n2684, B => n2579, Z => n2495);
   U2854 : ND2I port map( A => n2793, B => n2646, Z => n2679);
   U2855 : ND2I port map( A => n4835, B => n2702, Z => n2830);
   U2856 : ND2I port map( A => n2575, B => n2793, Z => n2702);
   U2859 : NR2I port map( A => n2582, B => n5054, Z => n1931);
   U2862 : ND2I port map( A => n2553, B => n2646, Z => n2515);
   U2864 : NR2I port map( A => n5075, B => n5060, Z => n2837);
   U2867 : NR2I port map( A => n2842, B => n2843, Z => n2841);
   U2869 : NR2I port map( A => n5045, B => n5061, Z => n2749);
   U2872 : AO1P port map( A => n5231, B => n2550, C => n2846, D => n2847, Z => 
                           n2840);
   U2875 : ND2I port map( A => n2668, B => n2657, Z => n2849);
   U2876 : NR2I port map( A => n5063, B => n5078, Z => n2848);
   U2878 : ND2I port map( A => n2521, B => n2793, Z => n2550);
   U2879 : ND2I port map( A => n5075, B => v_RAM_OUT0_24_port, Z => n2793);
   U2882 : ND2I port map( A => n2521, B => n4724, Z => n2855);
   U2883 : NR2I port map( A => n5076, B => n5054, Z => n2854);
   U2885 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2542, Z => n2574);
   U2887 : ND2I port map( A => n2732, B => n2707, Z => n2845);
   U2888 : ND2I port map( A => n2542, B => n4374, Z => n2707);
   U2889 : NR2I port map( A => n4828, B => n4510, Z => n2519);
   U2890 : ND2I port map( A => n2708, B => n2628, Z => n2856);
   U2891 : ND2I port map( A => n5078, B => n4374, Z => n2628);
   U2893 : ND2I port map( A => n2684, B => n2597, Z => n2670);
   U2897 : ND2I port map( A => n2860, B => n4432, Z => n2859);
   U2901 : ND2I port map( A => n4732, B => n4852, Z => n2483);
   U2902 : ND2I port map( A => n4852, B => n1674, Z => n2487);
   U2908 : ND2I port map( A => n4510, B => n4379, Z => n1924);
   U2913 : ND2I port map( A => n4835, B => n2714, Z => n2867);
   U2914 : ND2I port map( A => n2617, B => n2646, Z => n2714);
   U2915 : ND2I port map( A => n5074, B => n4374, Z => n2646);
   U2919 : ND2I port map( A => n2553, B => n2684, Z => n2642);
   U2920 : ND2I port map( A => v_RAM_OUT0_24_port, B => n4532, Z => n2553);
   U2921 : ND2I port map( A => n4724, B => n2542, Z => n1964);
   U2922 : ND2I port map( A => n2609, B => n2597, Z => n1962);
   U2923 : ND2I port map( A => n5076, B => v_RAM_OUT0_24_port, Z => n2597);
   U2925 : ND2I port map( A => v_RAM_OUT0_25_port, B => n4379, Z => n1922);
   U2928 : ND2I port map( A => n2752, B => n4724, Z => n2612);
   U2931 : NR2I port map( A => n5044, B => n5056, Z => n2647);
   U2933 : ND2I port map( A => v_RAM_OUT0_24_port, B => v_RAM_OUT0_27_port, Z 
                           => n2617);
   U2935 : ND2I port map( A => n4374, B => n2657, Z => n2534);
   U2937 : NR2I port map( A => n2618, B => n4397, Z => n2869);
   U2938 : ND2I port map( A => n5076, B => n4374, Z => n2618);
   U2940 : ND2I port map( A => n2609, B => n2579, Z => n2544);
   U2941 : ND2I port map( A => n5077, B => v_RAM_OUT0_24_port, Z => n2579);
   U2943 : ND2I port map( A => v_RAM_OUT0_30_port, B => n4416, Z => n2542);
   U2945 : ND2I port map( A => n4836, B => n4510, Z => n2577);
   U2946 : ND2I port map( A => n5060, B => n5233, Z => n2874);
   U2950 : NR2I port map( A => n5044, B => n5058, Z => n2583);
   U2952 : ND2I port map( A => n4532, B => n4374, Z => n2731);
   U2958 : ND2I port map( A => v_RAM_OUT0_29_port, B => n4510, Z => n2533);
   U2961 : NR2I port map( A => n5045, B => n5059, Z => n2645);
   U2964 : ND2I port map( A => n4374, B => n2752, Z => n2520);
   U2967 : ND2I port map( A => n5078, B => v_RAM_OUT0_24_port, Z => n1930);
   U2970 : ND2I port map( A => n4416, B => n4374, Z => n2521);
   U2973 : NR2I port map( A => n5058, B => n5047, Z => n1953);
   U2975 : ND2I port map( A => n5075, B => n4374, Z => n2516);
   U2978 : ND2I port map( A => n5074, B => v_RAM_OUT0_24_port, Z => n2708);
   U2980 : ND2I port map( A => n2499, B => n2684, Z => n2532);
   U2981 : ND2I port map( A => n2582, B => n4374, Z => n2684);
   U2982 : ND2I port map( A => v_RAM_OUT0_24_port, B => n4416, Z => n2499);
   U2984 : ND2I port map( A => n4725, B => n4828, Z => n1954);
   U2986 : ND2I port map( A => v_RAM_OUT0_25_port, B => v_RAM_OUT0_29_port, Z 
                           => n2536);
   U2989 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2582, Z => n2610);
   U2990 : ND2I port map( A => n2657, B => n2752, Z => n2582);
   U2991 : NR2I port map( A => n4727, B => v_RAM_OUT0_25_port, Z => n2524);
   U2993 : ND2I port map( A => n5234, B => n4510, Z => n2511);
   U2996 : ND2I port map( A => n2668, B => n2609, Z => n2801);
   U2997 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2752, Z => n2668);
   U2998 : ND2I port map( A => v_RAM_OUT0_27_port, B => v_RAM_OUT0_30_port, Z 
                           => n2752);
   U3000 : ND2I port map( A => n5231, B => v_RAM_OUT0_25_port, Z => n2526);
   U3002 : ND2I port map( A => n4781, B => n4397, Z => n1966);
   U3004 : ND2I port map( A => n5234, B => v_RAM_OUT0_25_port, Z => n2522);
   U3006 : ND2I port map( A => v_RAM_OUT0_26_port, B => n4781, Z => n2611);
   U3008 : ND2I port map( A => v_RAM_OUT0_24_port, B => v_RAM_OUT0_30_port, Z 
                           => n2732);
   U3009 : ND2I port map( A => n4834, B => n2721, Z => n2885);
   U3010 : ND2I port map( A => n4724, B => n2796, Z => n2721);
   U3011 : ND2I port map( A => n2575, B => n4374, Z => n2796);
   U3012 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2657, Z => n1949);
   U3013 : ND2I port map( A => n4532, B => n4416, Z => n2657);
   U3018 : ND2I port map( A => n2541, B => n2609, Z => n2815);
   U3021 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2575, Z => n2541);
   U3025 : ND2I port map( A => n4839, B => v_RAM_OUT0_25_port, Z => n2578);
   U3028 : ND2I port map( A => n4839, B => n4510, Z => n2644);
   U3031 : ND2I port map( A => v_RAM_OUT0_26_port, B => n4360, Z => n1929);
   U3036 : ND2I port map( A => n2891, B => n4534, Z => n2889);
   U3051 : NR2I port map( A => n4395, B => n4509, Z => n2925);
   U3060 : AO1P port map( A => n5194, B => n5087, C => n2947, D => n2948, Z => 
                           n2938);
   U3068 : ND2I port map( A => n2930, B => n2961, Z => n2908);
   U3075 : ND2I port map( A => n2969, B => n4423, Z => n2967);
   U3081 : AO1P port map( A => n2978, B => n4509, C => n2979, D => n2980, Z => 
                           n2977);
   U3084 : ND2I port map( A => n5093, B => n2988, Z => n2978);
   U3090 : ND2I port map( A => n5090, B => n4395, Z => n2998);
   U3093 : ND2I port map( A => n3004, B => n3005, Z => n2960);
   U3095 : ND2I port map( A => n3008, B => n3009, Z => n2971);
   U3097 : AO1P port map( A => n5220, B => n5097, C => n3013, D => n3014, Z => 
                           n3010);
   U3098 : NR2I port map( A => n4813, B => n2982, Z => n3014);
   U3101 : AO1P port map( A => n4817, B => n3020, C => n3021, D => n3022, Z => 
                           n3019);
   U3103 : NR2I port map( A => n5100, B => n4717, Z => n3021);
   U3109 : AO1P port map( A => n5223, B => n3032, C => n3033, D => n3034, Z => 
                           n3026);
   U3112 : ND2I port map( A => n3024, B => n3003, Z => n3032);
   U3116 : ND2I port map( A => n3038, B => n4422, Z => n3036);
   U3121 : NR2I port map( A => n3043, B => n3044, Z => n3042);
   U3130 : AO1P port map( A => n4817, B => n2958, C => v_RAM_OUT0_17_port, D =>
                           n3062, Z => n3061);
   U3131 : NR2I port map( A => n4718, B => n3015, Z => n3062);
   U3135 : NR2I port map( A => n4780, B => n5109, Z => n3067);
   U3136 : ND2I port map( A => v_RAM_OUT0_23_port, B => n3070, Z => n3041);
   U3138 : AO1P port map( A => n5220, B => n3073, C => n3074, D => n3075, Z => 
                           n3072);
   U3141 : ND2I port map( A => n2981, B => n2943, Z => n3073);
   U3151 : AO1P port map( A => n5112, B => n5220, C => n3093, D => n3094, Z => 
                           n3079);
   U3153 : NR2I port map( A => n5236, B => n5112, Z => n2964);
   U3157 : ND2I port map( A => n3099, B => n4553, Z => n3097);
   U3160 : ND2I port map( A => n3100, B => n3101, Z => n1628);
   U3169 : ND2I port map( A => n2943, B => n3114, Z => n3085);
   U3170 : NR2I port map( A => n5079, B => n5099, Z => n3091);
   U3172 : NR2I port map( A => n4782, B => n4813, Z => n3110);
   U3176 : ND2I port map( A => n3065, B => n3016, Z => n3107);
   U3180 : NR2I port map( A => n3120, B => n4717, Z => n3094);
   U3186 : NR2I port map( A => n5107, B => n5096, Z => n3128);
   U3193 : AO1P port map( A => n5220, B => n3134, C => n3135, D => n3136, Z => 
                           n3133);
   U3196 : ND2I port map( A => n2943, B => n2961, Z => n3134);
   U3203 : ND2I port map( A => n3145, B => n4614, Z => n3142);
   U3209 : ND2I port map( A => n3153, B => n3154, Z => n3152);
   U3214 : ND2I port map( A => n5223, B => n3065, Z => n3157);
   U3217 : ND2I port map( A => n5100, B => n2949, Z => n2966);
   U3221 : ND2I port map( A => n2930, B => n3138, Z => n3165);
   U3223 : ND2I port map( A => n3015, B => n3114, Z => n3168);
   U3224 : NR2I port map( A => n5097, B => n5114, Z => n3167);
   U3225 : NR2I port map( A => n5114, B => n5108, Z => n3162);
   U3228 : AO1P port map( A => n4815, B => n3090, C => n3173, D => n3174, Z => 
                           n3172);
   U3229 : NR2I port map( A => n4718, B => n3016, Z => n3174);
   U3231 : ND2I port map( A => n2906, B => n2924, Z => n3090);
   U3232 : AO1P port map( A => n5238, B => n5223, C => n3176, D => n3177, Z => 
                           n3171);
   U3235 : NR2I port map( A => n5090, B => n5239, Z => n2999);
   U3237 : AO1P port map( A => n5113, B => n5221, C => n3181, D => n3182, Z => 
                           n3179);
   U3238 : NR2I port map( A => n5114, B => n3183, Z => n3182);
   U3240 : AO1P port map( A => n4812, B => n3184, C => n1682, D => n4509, Z => 
                           n3181);
   U3241 : ND2I port map( A => n3185, B => n4395, Z => n3184);
   U3243 : ND2I port map( A => n3137, B => n3016, Z => n3185);
   U3247 : ND2I port map( A => n3189, B => n4613, Z => n3186);
   U3253 : AO1P port map( A => n5100, B => n1656, C => n3193, D => n3194, Z => 
                           n3192);
   U3254 : NR2I port map( A => n4823, B => n3003, Z => n3194);
   U3256 : ND2I port map( A => n3015, B => n3003, Z => n2932);
   U3263 : ND2I port map( A => n4819, B => n2982, Z => n3196);
   U3266 : ND2I port map( A => n4719, B => n3077, Z => n3202);
   U3268 : ND2I port map( A => n3024, B => n3016, Z => n3020);
   U3269 : AN2I port map( A => n3092, B => n3203, Z => n3108);
   U3277 : ND2I port map( A => n2930, B => n3076, Z => n3161);
   U3283 : ND2I port map( A => n2906, B => n3005, Z => n3215);
   U3284 : ND2I port map( A => n5108, B => n4373, Z => n3005);
   U3286 : ND2I port map( A => n3216, B => n3004, Z => n2991);
   U3287 : NR2I port map( A => n5110, B => n5238, Z => n3155);
   U3289 : ND2I port map( A => n4782, B => n4509, Z => n2942);
   U3292 : ND2I port map( A => n2986, B => n3113, Z => n2935);
   U3294 : ND2I port map( A => v_RAM_OUT0_17_port, B => n4782, Z => n2945);
   U3295 : NR2I port map( A => n3220, B => n3221, Z => n3207);
   U3298 : ND2I port map( A => n3159, B => n2981, Z => n3057);
   U3299 : NR2I port map( A => n5088, B => n5238, Z => n3141);
   U3301 : ND2I port map( A => v_RAM_OUT0_19_port, B => n4373, Z => n3077);
   U3305 : ND2I port map( A => n3225, B => n4561, Z => n3223);
   U3313 : ND2I port map( A => n2906, B => n3035, Z => n3007);
   U3319 : ND2I port map( A => n3092, B => n2986, Z => n2902);
   U3320 : ND2I port map( A => n3203, B => n3053, Z => n3087);
   U3321 : ND2I port map( A => n4820, B => n3109, Z => n3235);
   U3322 : ND2I port map( A => n2982, B => n3203, Z => n3109);
   U3326 : NR2I port map( A => n1657, B => n5110, Z => n1658);
   U3329 : ND2I port map( A => n2961, B => n3053, Z => n2922);
   U3331 : NR2I port map( A => n5100, B => n5114, Z => n3242);
   U3334 : NR2I port map( A => n3247, B => n3248, Z => n3246);
   U3336 : NR2I port map( A => n5115, B => n5105, Z => n3156);
   U3339 : AO1P port map( A => n5220, B => n2958, C => n3251, D => n3252, Z => 
                           n3245);
   U3342 : ND2I port map( A => n3076, B => n3065, Z => n3254);
   U3343 : NR2I port map( A => n5088, B => n5113, Z => n3253);
   U3345 : ND2I port map( A => n2930, B => n3203, Z => n2958);
   U3346 : ND2I port map( A => n5100, B => v_RAM_OUT0_16_port, Z => n3203);
   U3349 : ND2I port map( A => n2930, B => n4719, Z => n3260);
   U3350 : NR2I port map( A => n5087, B => n5110, Z => n3259);
   U3352 : ND2I port map( A => v_RAM_OUT0_16_port, B => n2950, Z => n2981);
   U3354 : ND2I port map( A => n3138, B => n3113, Z => n3250);
   U3355 : ND2I port map( A => n2950, B => n4373, Z => n3113);
   U3356 : NR2I port map( A => n4813, B => n4509, Z => n2927);
   U3357 : ND2I port map( A => n3114, B => n3035, Z => n3261);
   U3358 : ND2I port map( A => n5113, B => n4373, Z => n3035);
   U3360 : ND2I port map( A => n3092, B => n3004, Z => n3078);
   U3366 : ND2I port map( A => n3264, B => n4549, Z => n3262);
   U3369 : ND2I port map( A => n4722, B => n4852, Z => n2888);
   U3370 : ND2I port map( A => n4852, B => n1726, Z => n2892);
   U3377 : ND2I port map( A => n3076, B => n3015, Z => n3222);
   U3379 : ND2I port map( A => v_RAM_OUT0_16_port, B => v_RAM_OUT0_22_port, Z 
                           => n3138);
   U3380 : ND2I port map( A => n4820, B => n3127, Z => n3270);
   U3381 : ND2I port map( A => n4719, B => n3216, Z => n3127);
   U3382 : ND2I port map( A => n2982, B => n4373, Z => n3216);
   U3384 : ND2I port map( A => n2949, B => n3015, Z => n3204);
   U3385 : ND2I port map( A => v_RAM_OUT0_16_port, B => n2982, Z => n2949);
   U3386 : AO1P port map( A => n5224, B => n4719, C => n3273, D => n3274, Z => 
                           n3268);
   U3387 : AN2I port map( A => n5219, B => n1697, Z => n3274);
   U3388 : NR2I port map( A => n5096, B => n5099, Z => n1697);
   U3390 : ND2I port map( A => n5100, B => n4373, Z => n2924);
   U3393 : ND2I port map( A => n4356, B => v_RAM_OUT0_17_port, Z => n2985);
   U3397 : NR2I port map( A => n5115, B => n5237, Z => n3052);
   U3400 : ND2I port map( A => n4373, B => n3159, Z => n2928);
   U3403 : ND2I port map( A => n5113, B => v_RAM_OUT0_16_port, Z => n3003);
   U3406 : ND2I port map( A => n4399, B => n4373, Z => n2930);
   U3410 : ND2I port map( A => v_RAM_OUT0_17_port, B => n4403, Z => n2901);
   U3414 : ND2I port map( A => n2961, B => n3092, Z => n3049);
   U3415 : ND2I port map( A => v_RAM_OUT0_16_port, B => n4512, Z => n2961);
   U3416 : ND2I port map( A => n4719, B => n2950, Z => n1685);
   U3417 : ND2I port map( A => n3015, B => n3004, Z => n1682);
   U3418 : ND2I port map( A => n5087, B => v_RAM_OUT0_16_port, Z => n3004);
   U3419 : ND2I port map( A => n4717, B => n4813, Z => n1684);
   U3420 : ND2I port map( A => n4509, B => n4402, Z => n2899);
   U3426 : ND2I port map( A => n2906, B => n3092, Z => n1694);
   U3427 : ND2I port map( A => n1657, B => n4373, Z => n3092);
   U3428 : ND2I port map( A => v_RAM_OUT0_16_port, B => n4399, Z => n2906);
   U3429 : ND2I port map( A => n4821, B => n3120, Z => n3282);
   U3430 : ND2I port map( A => n3023, B => n3053, Z => n3120);
   U3431 : ND2I port map( A => n5097, B => n4373, Z => n3053);
   U3434 : ND2I port map( A => n5223, B => n4509, Z => n2918);
   U3435 : ND2I port map( A => n3159, B => n4719, Z => n3018);
   U3436 : ND2I port map( A => v_RAM_OUT0_16_port, B => n3065, Z => n1696);
   U3439 : NR2I port map( A => n5104, B => n5239, Z => n3055);
   U3441 : ND2I port map( A => v_RAM_OUT0_16_port, B => v_RAM_OUT0_19_port, Z 
                           => n3023);
   U3443 : ND2I port map( A => n4373, B => n3065, Z => n2943);
   U3445 : NR2I port map( A => n3024, B => n4395, Z => n3284);
   U3446 : ND2I port map( A => n5087, B => n4373, Z => n3024);
   U3450 : ND2I port map( A => n3015, B => n2986, Z => n2951);
   U3451 : ND2I port map( A => n5108, B => v_RAM_OUT0_16_port, Z => n2986);
   U3453 : ND2I port map( A => v_RAM_OUT0_22_port, B => n4399, Z => n2950);
   U3456 : ND2I port map( A => n4819, B => n4509, Z => n2984);
   U3459 : ND2I port map( A => v_RAM_OUT0_16_port, B => n1657, Z => n3016);
   U3461 : ND2I port map( A => n5220, B => v_RAM_OUT0_17_port, Z => n2936);
   U3463 : ND2I port map( A => n5114, B => n5222, Z => n3286);
   U3465 : ND2I port map( A => n5223, B => v_RAM_OUT0_17_port, Z => n2931);
   U3467 : ND2I port map( A => v_RAM_OUT0_18_port, B => n4780, Z => n3017);
   U3469 : ND2I port map( A => v_RAM_OUT0_16_port, B => n3159, Z => n3076);
   U3472 : ND2I port map( A => n3065, B => n3159, Z => n1657);
   U3473 : ND2I port map( A => v_RAM_OUT0_19_port, B => v_RAM_OUT0_22_port, Z 
                           => n3159);
   U3475 : ND2I port map( A => n4356, B => n4509, Z => n3051);
   U3481 : NR2I port map( A => n5104, B => n5096, Z => n2989);
   U3483 : ND2I port map( A => n5097, B => v_RAM_OUT0_16_port, Z => n3114);
   U3485 : ND2I port map( A => n4512, B => n4399, Z => n3065);
   U3488 : ND2I port map( A => n4512, B => n4373, Z => n3137);
   U3491 : NR2I port map( A => n4714, B => v_RAM_OUT0_17_port, Z => n2934);
   U3492 : ND2I port map( A => n4780, B => n4395, Z => n2905);
   U3497 : ND2I port map( A => n3294, B => n4431, Z => n3292);
   U3511 : NR2I port map( A => n4371, B => n4508, Z => n3328);
   U3520 : AO1P port map( A => n5207, B => n5164, C => n3350, D => n3351, Z => 
                           n3341);
   U3528 : ND2I port map( A => n3333, B => n3364, Z => n3311);
   U3535 : ND2I port map( A => n3372, B => n4406, Z => n3370);
   U3540 : AO1P port map( A => n3381, B => n4508, C => n3382, D => n3383, Z => 
                           n3380);
   U3543 : ND2I port map( A => n5170, B => n3391, Z => n3381);
   U3549 : ND2I port map( A => n5167, B => n4371, Z => n3401);
   U3552 : ND2I port map( A => n3407, B => n3408, Z => n3363);
   U3554 : ND2I port map( A => n3411, B => n3412, Z => n3374);
   U3556 : AO1P port map( A => n5211, B => n5174, C => n3416, D => n3417, Z => 
                           n3413);
   U3557 : NR2I port map( A => n4797, B => n3385, Z => n3417);
   U3560 : AO1P port map( A => n4801, B => n3423, C => n3424, D => n3425, Z => 
                           n3422);
   U3562 : NR2I port map( A => n5177, B => n4707, Z => n3424);
   U3568 : AO1P port map( A => n5214, B => n3435, C => n3436, D => n3437, Z => 
                           n3429);
   U3571 : ND2I port map( A => n3427, B => n3406, Z => n3435);
   U3575 : ND2I port map( A => n3441, B => n4523, Z => n3439);
   U3579 : NR2I port map( A => n3446, B => n3447, Z => n3445);
   U3588 : AO1P port map( A => n4801, B => n3361, C => v_RAM_OUT0_1_port, D => 
                           n3465, Z => n3464);
   U3589 : NR2I port map( A => n4708, B => n3418, Z => n3465);
   U3593 : NR2I port map( A => n4779, B => n5186, Z => n3470);
   U3594 : ND2I port map( A => v_RAM_OUT0_7_port, B => n3473, Z => n3444);
   U3596 : AO1P port map( A => n5211, B => n3476, C => n3477, D => n3478, Z => 
                           n3475);
   U3599 : ND2I port map( A => n3384, B => n3346, Z => n3476);
   U3609 : AO1P port map( A => n5189, B => n5211, C => n3496, D => n3497, Z => 
                           n3482);
   U3611 : NR2I port map( A => n5243, B => n5189, Z => n3367);
   U3615 : ND2I port map( A => n3503, B => n4609, Z => n3500);
   U3617 : ND2I port map( A => n3504, B => n3505, Z => n1539);
   U3626 : ND2I port map( A => n3346, B => n3518, Z => n3488);
   U3627 : NR2I port map( A => n5156, B => n5176, Z => n3494);
   U3629 : NR2I port map( A => v_RAM_OUT0_5_port, B => n4797, Z => n3514);
   U3633 : ND2I port map( A => n3468, B => n3419, Z => n3511);
   U3637 : NR2I port map( A => n3524, B => n4707, Z => n3497);
   U3643 : NR2I port map( A => n5184, B => n5173, Z => n3532);
   U3650 : AO1P port map( A => n5211, B => n3538, C => n3539, D => n3540, Z => 
                           n3537);
   U3653 : ND2I port map( A => n3346, B => n3364, Z => n3538);
   U3660 : ND2I port map( A => n3549, B => n4608, Z => n3546);
   U3665 : ND2I port map( A => n3557, B => n3558, Z => n3556);
   U3670 : ND2I port map( A => n5214, B => n3468, Z => n3561);
   U3673 : ND2I port map( A => n5177, B => n3352, Z => n3369);
   U3677 : ND2I port map( A => n3333, B => n3542, Z => n3569);
   U3679 : ND2I port map( A => n3418, B => n3518, Z => n3572);
   U3680 : NR2I port map( A => n5174, B => n5191, Z => n3571);
   U3681 : NR2I port map( A => n5191, B => n5185, Z => n3566);
   U3684 : AO1P port map( A => n4799, B => n3493, C => n3577, D => n3578, Z => 
                           n3576);
   U3685 : NR2I port map( A => n4708, B => n3419, Z => n3578);
   U3687 : ND2I port map( A => n3309, B => n3327, Z => n3493);
   U3688 : AO1P port map( A => n5245, B => n5214, C => n3580, D => n3581, Z => 
                           n3575);
   U3691 : NR2I port map( A => n5167, B => n5246, Z => n3402);
   U3693 : AO1P port map( A => n5190, B => n5212, C => n3585, D => n3586, Z => 
                           n3583);
   U3694 : NR2I port map( A => n5191, B => n3587, Z => n3586);
   U3696 : AO1P port map( A => n4796, B => n3588, C => n2467, D => n4508, Z => 
                           n3585);
   U3697 : ND2I port map( A => n3589, B => n4371, Z => n3588);
   U3699 : ND2I port map( A => n3541, B => n3419, Z => n3589);
   U3703 : ND2I port map( A => n3593, B => n4607, Z => n3590);
   U3708 : AO1P port map( A => n5177, B => n2445, C => n3597, D => n3598, Z => 
                           n3596);
   U3709 : NR2I port map( A => n4807, B => n3406, Z => n3598);
   U3711 : ND2I port map( A => n3418, B => n3406, Z => n3335);
   U3718 : ND2I port map( A => n4803, B => n3385, Z => n3600);
   U3721 : ND2I port map( A => n4709, B => n3480, Z => n3606);
   U3723 : ND2I port map( A => n3427, B => n3419, Z => n3423);
   U3724 : AN2I port map( A => n3495, B => n3607, Z => n3512);
   U3732 : ND2I port map( A => n3333, B => n3479, Z => n3565);
   U3738 : ND2I port map( A => n3309, B => n3408, Z => n3619);
   U3739 : ND2I port map( A => n5185, B => n4372, Z => n3408);
   U3741 : ND2I port map( A => n3620, B => n3407, Z => n3394);
   U3742 : NR2I port map( A => n5187, B => n5245, Z => n3559);
   U3744 : ND2I port map( A => v_RAM_OUT0_5_port, B => n4508, Z => n3345);
   U3747 : ND2I port map( A => n3389, B => n3517, Z => n3338);
   U3749 : ND2I port map( A => v_RAM_OUT0_1_port, B => v_RAM_OUT0_5_port, Z => 
                           n3348);
   U3750 : NR2I port map( A => n3624, B => n3625, Z => n3611);
   U3753 : ND2I port map( A => n3563, B => n3384, Z => n3460);
   U3754 : NR2I port map( A => n5165, B => n5245, Z => n3545);
   U3756 : ND2I port map( A => v_RAM_OUT0_3_port, B => n4372, Z => n3480);
   U3760 : ND2I port map( A => n3630, B => n4606, Z => n3627);
   U3767 : ND2I port map( A => n3309, B => n3438, Z => n3410);
   U3773 : ND2I port map( A => n3495, B => n3389, Z => n3305);
   U3774 : ND2I port map( A => n3607, B => n3456, Z => n3490);
   U3775 : ND2I port map( A => n4804, B => n3513, Z => n3640);
   U3776 : ND2I port map( A => n3385, B => n3607, Z => n3513);
   U3780 : NR2I port map( A => n2446, B => n5187, Z => n2447);
   U3783 : ND2I port map( A => n3364, B => n3456, Z => n3325);
   U3785 : NR2I port map( A => n5177, B => n5191, Z => n3647);
   U3788 : NR2I port map( A => n3652, B => n3653, Z => n3651);
   U3790 : NR2I port map( A => n5192, B => n5182, Z => n3560);
   U3793 : AO1P port map( A => n5211, B => n3361, C => n3656, D => n3657, Z => 
                           n3650);
   U3796 : ND2I port map( A => n3479, B => n3468, Z => n3659);
   U3797 : NR2I port map( A => n5165, B => n5190, Z => n3658);
   U3799 : ND2I port map( A => n3333, B => n3607, Z => n3361);
   U3800 : ND2I port map( A => n5177, B => v_RAM_OUT0_0_port, Z => n3607);
   U3803 : ND2I port map( A => n3333, B => n4709, Z => n3665);
   U3804 : NR2I port map( A => n5164, B => n5187, Z => n3664);
   U3806 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3353, Z => n3384);
   U3808 : ND2I port map( A => n3542, B => n3517, Z => n3655);
   U3809 : ND2I port map( A => n3353, B => n4372, Z => n3517);
   U3810 : NR2I port map( A => n4797, B => n4508, Z => n3330);
   U3811 : ND2I port map( A => n3518, B => n3438, Z => n3666);
   U3812 : ND2I port map( A => n5190, B => n4372, Z => n3438);
   U3814 : ND2I port map( A => n3495, B => n3407, Z => n3481);
   U3820 : ND2I port map( A => n3670, B => n4605, Z => n3667);
   U3822 : ND2I port map( A => n4712, B => n4856, Z => n3291);
   U3823 : ND2I port map( A => n4857, B => n1726, Z => n3295);
   U3824 : ND2I port map( A => n3671, B => n4556, Z => n1726);
   U3833 : ND2I port map( A => n3479, B => n3418, Z => n3626);
   U3835 : ND2I port map( A => v_RAM_OUT0_0_port, B => v_RAM_OUT0_6_port, Z => 
                           n3542);
   U3836 : ND2I port map( A => n4804, B => n3531, Z => n3678);
   U3837 : ND2I port map( A => n4709, B => n3620, Z => n3531);
   U3838 : ND2I port map( A => n3385, B => n4372, Z => n3620);
   U3840 : ND2I port map( A => n3352, B => n3418, Z => n3608);
   U3841 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3385, Z => n3352);
   U3842 : AO1P port map( A => n5215, B => n4709, C => n3681, D => n3682, Z => 
                           n3676);
   U3843 : AN2I port map( A => n5210, B => n2482, Z => n3682);
   U3844 : NR2I port map( A => n5173, B => n5176, Z => n2482);
   U3846 : ND2I port map( A => n5177, B => n4372, Z => n3327);
   U3849 : ND2I port map( A => n4808, B => v_RAM_OUT0_1_port, Z => n3388);
   U3853 : NR2I port map( A => n5192, B => n5244, Z => n3455);
   U3856 : ND2I port map( A => n4372, B => n3563, Z => n3331);
   U3859 : ND2I port map( A => n5190, B => v_RAM_OUT0_0_port, Z => n3406);
   U3862 : ND2I port map( A => n4398, B => n4372, Z => n3333);
   U3866 : ND2I port map( A => v_RAM_OUT0_1_port, B => n4401, Z => n3304);
   U3870 : ND2I port map( A => n3364, B => n3495, Z => n3452);
   U3871 : ND2I port map( A => v_RAM_OUT0_0_port, B => n4511, Z => n3364);
   U3872 : ND2I port map( A => n4709, B => n3353, Z => n2470);
   U3873 : ND2I port map( A => n3418, B => n3407, Z => n2467);
   U3874 : ND2I port map( A => n5164, B => v_RAM_OUT0_0_port, Z => n3407);
   U3875 : ND2I port map( A => n4707, B => n4797, Z => n2469);
   U3876 : ND2I port map( A => n4508, B => n4401, Z => n3302);
   U3882 : ND2I port map( A => n3309, B => n3495, Z => n2479);
   U3883 : ND2I port map( A => n2446, B => n4372, Z => n3495);
   U3884 : ND2I port map( A => v_RAM_OUT0_0_port, B => n4398, Z => n3309);
   U3885 : ND2I port map( A => n4805, B => n3524, Z => n3690);
   U3886 : ND2I port map( A => n3426, B => n3456, Z => n3524);
   U3887 : ND2I port map( A => n5174, B => n4372, Z => n3456);
   U3890 : ND2I port map( A => n5214, B => n4508, Z => n3321);
   U3891 : ND2I port map( A => n3563, B => n4709, Z => n3421);
   U3892 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3468, Z => n2481);
   U3895 : NR2I port map( A => n5181, B => n5246, Z => n3458);
   U3897 : ND2I port map( A => v_RAM_OUT0_0_port, B => v_RAM_OUT0_3_port, Z => 
                           n3426);
   U3899 : ND2I port map( A => n4372, B => n3468, Z => n3346);
   U3901 : NR2I port map( A => n3427, B => n4371, Z => n3692);
   U3902 : ND2I port map( A => n5164, B => n4372, Z => n3427);
   U3906 : ND2I port map( A => n3418, B => n3389, Z => n3354);
   U3907 : ND2I port map( A => n5185, B => v_RAM_OUT0_0_port, Z => n3389);
   U3909 : ND2I port map( A => v_RAM_OUT0_6_port, B => n4398, Z => n3353);
   U3912 : ND2I port map( A => n4803, B => n4508, Z => n3387);
   U3915 : ND2I port map( A => v_RAM_OUT0_0_port, B => n2446, Z => n3419);
   U3917 : ND2I port map( A => n5211, B => v_RAM_OUT0_1_port, Z => n3339);
   U3919 : ND2I port map( A => n5191, B => n5213, Z => n3694);
   U3921 : ND2I port map( A => n5214, B => v_RAM_OUT0_1_port, Z => n3334);
   U3923 : ND2I port map( A => v_RAM_OUT0_2_port, B => n4779, Z => n3420);
   U3925 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3563, Z => n3479);
   U3928 : ND2I port map( A => n3468, B => n3563, Z => n2446);
   U3929 : ND2I port map( A => v_RAM_OUT0_3_port, B => v_RAM_OUT0_6_port, Z => 
                           n3563);
   U3931 : ND2I port map( A => n4808, B => n4508, Z => n3454);
   U3934 : ND2I port map( A => v_RAM_OUT0_2_port, B => n4358, Z => n3310);
   U3937 : NR2I port map( A => n5181, B => n5173, Z => n3392);
   U3939 : ND2I port map( A => n5174, B => v_RAM_OUT0_0_port, Z => n3518);
   U3941 : ND2I port map( A => n4511, B => n4398, Z => n3468);
   U3944 : ND2I port map( A => n4511, B => n4372, Z => n3541);
   U3947 : NR2I port map( A => n4704, B => v_RAM_OUT0_1_port, Z => n3337);
   U3948 : ND2I port map( A => n4779, B => n4371, Z => n3308);
   U3951 : ND2I port map( A => n4703, B => n3699, Z => N192);
   U3953 : ND2I port map( A => n1386, B => n4380, Z => n1388);
   U3955 : NR2I port map( A => n4540, B => n4999, Z => n1386);
   U3957 : ND2I port map( A => n3700, B => n3701, Z => n4314);
   U3961 : ND2I port map( A => n3954, B => n1433, Z => n1440);
   U3965 : ND2I port map( A => CE_I, B => n5010, Z => n3704);
   U3973 : AO1P port map( A => n4700, B => n4546, C => n3716, D => n3717, Z => 
                           n3715);
   U3995 : AO1P port map( A => n4700, B => n4430, C => n3729, D => n3730, Z => 
                           n3728);
   U4017 : AO1P port map( A => n4700, B => n4528, C => n3741, D => n3742, Z => 
                           n3740);
   U4039 : AO1P port map( A => n4700, B => n4583, C => n3752, D => n3753, Z => 
                           n3751);
   U4061 : AO1P port map( A => n4700, B => n4451, C => n3763, D => n3764, Z => 
                           n3762);
   U4083 : AO1P port map( A => n4700, B => n4582, C => n3774, D => n3775, Z => 
                           n3773);
   U4105 : AO1P port map( A => n4700, B => n4581, C => n3785, D => n3786, Z => 
                           n3784);
   U4125 : ND2I port map( A => n4353, B => n5016, Z => n1484);
   U4127 : ND2I port map( A => n1353, B => n4604, Z => n1343);
   U4131 : ND2I port map( A => n4352, B => n5021, Z => n1572);
   U4135 : AO1P port map( A => n4700, B => n4429, C => n3796, D => n3797, Z => 
                           n3795);
   U4138 : NR2I port map( A => n3798, B => n3799, Z => n1479);
   U4140 : NR2I port map( A => n5018, B => n3799, Z => n1478);
   U4145 : NR2I port map( A => n2376, B => n3802, Z => n1475);
   U4147 : NR2I port map( A => n3802, B => n2861, Z => n1476);
   U4149 : NR2I port map( A => n3799, B => n2376, Z => n1477);
   U4152 : ND2I port map( A => n3804, B => n3800, Z => n1469);
   U4153 : ND2I port map( A => n3800, B => n3805, Z => n1470);
   U4154 : NR2I port map( A => n4604, B => v_CALCULATION_CNTR_2_port, Z => 
                           n3800);
   U4156 : NR2I port map( A => n5024, B => n2861, Z => n1472);
   U4159 : NR2I port map( A => n3798, B => n5025, Z => n1467);
   U4161 : NR2I port map( A => n3799, B => n2861, Z => n1465);
   U4162 : ND2I port map( A => v_CALCULATION_CNTR_0_port, B => 
                           v_CALCULATION_CNTR_2_port, Z => n2861);
   U4163 : ND2I port map( A => v_CALCULATION_CNTR_3_port, B => n5026, Z => 
                           n3799);
   U4167 : NR2I port map( A => n5024, B => n3798, Z => n1473);
   U4168 : ND2I port map( A => n4556, B => n4604, Z => n3798);
   U4171 : NR2I port map( A => n5024, B => n2376, Z => n1466);
   U4175 : ND2I port map( A => n4411, B => n4369, Z => n2377);
   U4178 : ND2I port map( A => n1353, B => v_CALCULATION_CNTR_0_port, Z => 
                           n1444);
   U4179 : NR2I port map( A => n3802, B => v_CALCULATION_CNTR_2_port, Z => 
                           n1353);
   U4184 : ND2I port map( A => n4439, B => n3672, Z => n3708);
   U4185 : ND2I port map( A => v_CALCULATION_CNTR_2_port, B => n3671, Z => 
                           n3672);
   U4187 : ND2I port map( A => v_CALCULATION_CNTR_1_port, B => n1458, Z => 
                           n1457);
   U4188 : NR4P port map( A => v_CALCULATION_CNTR_4_port, B => 
                           v_CALCULATION_CNTR_5_port, C => 
                           v_CALCULATION_CNTR_6_port, D => 
                           v_CALCULATION_CNTR_7_port, Z => n1458);
   U4195 : NR2I port map( A => RESET_I, B => n3957, Z => n1433);
   U4197 : NR2I port map( A => n5025, B => n2376, Z => n1474);
   U4198 : ND2I port map( A => v_CALCULATION_CNTR_2_port, B => n4604, Z => 
                           n2376);
   U4205 : ND2I port map( A => n5010, B => n4892, Z => n1413);
   KEXP0 : key_expansion port map( KEY_I(7) => KEY_I(7), KEY_I(6) => KEY_I(6), 
                           KEY_I(5) => KEY_I(5), KEY_I(4) => KEY_I(4), KEY_I(3)
                           => KEY_I(3), KEY_I(2) => KEY_I(2), KEY_I(1) => 
                           KEY_I(1), KEY_I(0) => KEY_I(0), VALID_KEY_I => 
                           VALID_KEY_I, CLK_I => CLK_I, RESET_I => RESET_I, 
                           CE_I => CE_I, DONE_O => KEY_READY_O, GET_KEY_I => 
                           GET_KEY, KEY_NUMB_I(5) => v_INV_KEY_NUMB_5_port, 
                           KEY_NUMB_I(4) => v_INV_KEY_NUMB_4_port, 
                           KEY_NUMB_I(3) => v_INV_KEY_NUMB_3_port, 
                           KEY_NUMB_I(2) => v_INV_KEY_NUMB_2_port, 
                           KEY_NUMB_I(1) => n4666, KEY_NUMB_I(0) => n4667, 
                           KEY_EXP_O(31) => v_KEY_COLUMN_31_port, KEY_EXP_O(30)
                           => v_KEY_COLUMN_30_port, KEY_EXP_O(29) => 
                           v_KEY_COLUMN_29_port, KEY_EXP_O(28) => 
                           v_KEY_COLUMN_28_port, KEY_EXP_O(27) => 
                           v_KEY_COLUMN_27_port, KEY_EXP_O(26) => 
                           v_KEY_COLUMN_26_port, KEY_EXP_O(25) => 
                           v_KEY_COLUMN_25_port, KEY_EXP_O(24) => 
                           v_KEY_COLUMN_24_port, KEY_EXP_O(23) => 
                           v_KEY_COLUMN_23_port, KEY_EXP_O(22) => 
                           v_KEY_COLUMN_22_port, KEY_EXP_O(21) => 
                           v_KEY_COLUMN_21_port, KEY_EXP_O(20) => 
                           v_KEY_COLUMN_20_port, KEY_EXP_O(19) => 
                           v_KEY_COLUMN_19_port, KEY_EXP_O(18) => 
                           v_KEY_COLUMN_18_port, KEY_EXP_O(17) => 
                           v_KEY_COLUMN_17_port, KEY_EXP_O(16) => 
                           v_KEY_COLUMN_16_port, KEY_EXP_O(15) => 
                           v_KEY_COLUMN_15_port, KEY_EXP_O(14) => 
                           v_KEY_COLUMN_14_port, KEY_EXP_O(13) => 
                           v_KEY_COLUMN_13_port, KEY_EXP_O(12) => 
                           v_KEY_COLUMN_12_port, KEY_EXP_O(11) => 
                           v_KEY_COLUMN_11_port, KEY_EXP_O(10) => 
                           v_KEY_COLUMN_10_port, KEY_EXP_O(9) => 
                           v_KEY_COLUMN_9_port, KEY_EXP_O(8) => 
                           v_KEY_COLUMN_8_port, KEY_EXP_O(7) => 
                           v_KEY_COLUMN_7_port, KEY_EXP_O(6) => 
                           v_KEY_COLUMN_6_port, KEY_EXP_O(5) => 
                           v_KEY_COLUMN_5_port, KEY_EXP_O(4) => 
                           v_KEY_COLUMN_4_port, KEY_EXP_O(3) => 
                           v_KEY_COLUMN_3_port, KEY_EXP_O(2) => 
                           v_KEY_COLUMN_2_port, KEY_EXP_O(1) => 
                           v_KEY_COLUMN_1_port, KEY_EXP_O(0) => 
                           v_KEY_COLUMN_0_port);
   U4208 : AO2 port map( A => n4920, B => n196, C => n198, D => n1336, Z => 
                           n1335);
   U4209 : AO2 port map( A => n196, B => n1336, C => n4920, D => n198, Z => 
                           n1333);
   U4210 : NR2I port map( A => n1339, B => n1340, Z => n196);
   U4211 : AO3 port map( A => n4886, B => n4472, C => n1278, D => n1279, Z => 
                           n3974);
   U4212 : AO3 port map( A => n4886, B => n4473, C => n970, D => n971, Z => 
                           n3980);
   U4213 : AO3 port map( A => n4888, B => n4474, C => n145, D => n146, Z => 
                           n3986);
   U4214 : EON1 port map( A => n4411, B => n1413, C => N2083, D => n1409, Z => 
                           n4312);
   U4215 : AN2I port map( A => v_RAM_OUT0_18_port, B => n4355, Z => n4356);
   U4216 : ND2I port map( A => n3948, B => n1426, Z => n4361);
   U4217 : ND3 port map( A => n1424, B => n3949, C => n3948, Z => n4362);
   U4218 : NR3P port map( A => n4892, B => n3943, C => n4366, Z => n4363);
   U4219 : ND3 port map( A => n4603, B => n4366, C => CE_I, Z => n4367);
   U4220 : ND4P port map( A => n5023, B => n4886, C => n5015, D => n5010, Z => 
                           n4368);
   U4221 : AN3 port map( A => n1315, B => n4886, C => n5016, Z => n4370);
   U4222 : AN2I port map( A => n5023, B => n4439, Z => n4381);
   U4223 : AN2I port map( A => n1426, B => n4466, Z => n4393);
   U4224 : AN3 port map( A => n4466, B => n1424, C => n3949, Z => n4394);
   U4225 : AN2I port map( A => n4352, B => n5022, Z => n4396);
   U4226 : ND4 port map( A => n1315, B => n4886, C => n1342, D => n1343, Z => 
                           n1340);
   U4227 : AN2I port map( A => n4395, B => n4354, Z => n4505);
   U4228 : AN2I port map( A => n4371, B => n4357, Z => n4513);
   U4229 : AN2I port map( A => n4397, B => n4359, Z => n4514);
   U4230 : OR2P port map( A => n103, B => n3942, Z => n4584);
   U4231 : OR2P port map( A => n4366, B => n103, Z => n4585);
   U4232 : IVI port map( A => n4854, Z => n4852);
   U4233 : IVI port map( A => n4821, Z => n4813);
   U4234 : IVI port map( A => n4854, Z => n4850);
   U4235 : IVI port map( A => n4854, Z => n4849);
   U4236 : IVI port map( A => n4854, Z => n4851);
   U4237 : IVI port map( A => n4848, Z => n4845);
   U4238 : IVI port map( A => n4848, Z => n4846);
   U4239 : IVI port map( A => n4805, Z => n4797);
   U4240 : IVI port map( A => n4836, Z => n4828);
   U4241 : IVI port map( A => n4848, Z => n4843);
   U4242 : IVI port map( A => n4848, Z => n4844);
   U4243 : IVI port map( A => n4819, Z => n4812);
   U4244 : IVI port map( A => n4803, Z => n4796);
   U4245 : IVDA port map( A => n4506, Y => n4364, Z => n4767);
   U4246 : IVDA port map( A => n4506, Y => n4365, Z => n4768);
   U4247 : IVI port map( A => n4834, Z => n4827);
   U4248 : IVI port map( A => n4884, Z => n4865);
   U4249 : IVI port map( A => n4884, Z => n4866);
   U4250 : IVI port map( A => n4396, Z => n4842);
   U4251 : IVDA port map( A => n2001, Y => n_3395, Z => n4741);
   U4252 : IVDA port map( A => n1530, Y => n_3396, Z => n4759);
   U4253 : IVDA port map( A => n2001, Y => n_3397, Z => n4742);
   U4254 : AO2 port map( A => n5199, B => n5129, C => n5197, D => n5136, Z => 
                           n2026);
   U4255 : IVDA port map( A => n1530, Y => n_3398, Z => n4760);
   U4256 : IVI port map( A => n4396, Z => n4840);
   U4257 : IVI port map( A => n4396, Z => n4841);
   U4258 : IVDA port map( A => n4507, Y => n4376, Z => n4765);
   U4259 : IVDA port map( A => n4507, Y => n4377, Z => n4766);
   U4260 : IVDA port map( A => n4504, Y => n4413, Z => n4770);
   U4261 : IVDA port map( A => n1791, Y => n_3399, Z => n4749);
   U4262 : IVDA port map( A => n4515, Y => n4412, Z => n4769);
   U4263 : IVDA port map( A => n1791, Y => n_3400, Z => n4750);
   U4264 : AO2 port map( A => n1005, B => n196, C => n198, D => n4919, Z => 
                           n1003);
   U4265 : AO2 port map( A => n196, B => n4919, C => n1005, D => n198, Z => 
                           n1001);
   U4266 : AO2 port map( A => n4932, B => n196, C => n197, D => n198, Z => n193
                           );
   U4267 : AO2 port map( A => n197, B => n196, C => n4932, D => n198, Z => n191
                           );
   U4268 : AO4 port map( A => n1333, B => n4912, C => n1335, D => n655, Z => 
                           n1332);
   U4269 : AO4 port map( A => n1333, B => n655, C => n1335, D => n4912, Z => 
                           n1331);
   U4270 : IVI port map( A => n4370, Z => n4885);
   U4271 : IVI port map( A => n4792, Z => n4789);
   U4272 : IVI port map( A => n4786, Z => n4783);
   U4273 : IVI port map( A => n1340, Z => n4787);
   U4274 : IVI port map( A => n4792, Z => n4790);
   U4275 : IVI port map( A => n4786, Z => n4784);
   U4276 : IVI port map( A => n1340, Z => n4788);
   U4277 : AO4 port map( A => n4885, B => n336, C => n4368, D => n337, Z => 
                           n335);
   U4278 : AO4 port map( A => n4885, B => n667, C => n4368, D => n668, Z => 
                           n666);
   U4279 : IVDA port map( A => n1972, Y => n_3401, Z => n4743);
   U4280 : IVDA port map( A => n2414, Y => n_3402, Z => n4734);
   U4281 : EON1 port map( A => n5080, B => n2984, C => n3053, D => n5219, Z => 
                           n3046);
   U4282 : EON1 port map( A => n5157, B => n3387, C => n3456, D => n5210, Z => 
                           n3449);
   U4283 : IVDA port map( A => n1898, Y => n_3403, Z => n4745);
   U4284 : IVDA port map( A => n2487, Y => n_3404, Z => n4732);
   U4285 : IVDA port map( A => n2892, Y => n_3405, Z => n4722);
   U4286 : IVDA port map( A => n1898, Y => n_3406, Z => n4746);
   U4287 : IVDA port map( A => n1972, Y => n_3407, Z => n4744);
   U4288 : IVDA port map( A => n2414, Y => n_3408, Z => n4735);
   U4289 : IVI port map( A => n1474, Z => n5020);
   U4290 : AO2 port map( A => n2991, B => n5220, C => n5223, D => n5110, Z => 
                           n3060);
   U4291 : AO2 port map( A => n3394, B => n5211, C => n5214, D => n5187, Z => 
                           n3463);
   U4292 : AO4 port map( A => n4413, B => n2111, C => n2180, D => n4739, Z => 
                           n2179);
   U4293 : AO7 port map( A => n4736, B => n2035, C => n5070, Z => n2178);
   U4294 : IVI port map( A => n2210, Z => n5197);
   U4295 : IVI port map( A => n2076, Z => n5199);
   U4296 : EON1 port map( A => n2319, B => n4738, C => n2035, D => n4504, Z => 
                           n2366);
   U4297 : AO7 port map( A => n1888, B => n5235, C => n2390, Z => n2385);
   U4298 : AO2 port map( A => n1890, B => n4504, C => n4507, D => n1889, Z => 
                           n2390);
   U4299 : AO2 port map( A => n5198, B => n5135, C => n1888, D => n5196, Z => 
                           n2368);
   U4300 : AO2 port map( A => n5201, B => n1884, C => n5143, D => n5203, Z => 
                           n2171);
   U4301 : IVDA port map( A => n1617, Y => n_3409, Z => n4757);
   U4302 : IVDA port map( A => n1702, Y => n_3410, Z => n4755);
   U4303 : IVDA port map( A => n1731, Y => n_3411, Z => n4753);
   U4304 : IVDA port map( A => n2487, Y => n_3412, Z => n4733);
   U4305 : IVDA port map( A => n2892, Y => n_3413, Z => n4723);
   U4306 : IVDA port map( A => n1617, Y => n_3414, Z => n4758);
   U4307 : IVDA port map( A => n1702, Y => n_3415, Z => n4756);
   U4308 : IVDA port map( A => n1731, Y => n_3416, Z => n4754);
   U4309 : AO2 port map( A => n2585, B => n5231, C => n5234, D => n5054, Z => 
                           n2652);
   U4310 : IVI port map( A => n2070, Z => n5198);
   U4311 : NR3 port map( A => n4738, B => n5134, C => n5130, Z => n2101);
   U4312 : IVI port map( A => n2078, Z => n5196);
   U4313 : AO7 port map( A => n5053, B => n5044, C => n4839, Z => n2791);
   U4314 : AO7 port map( A => n5098, B => n5104, C => n4356, Z => n3212);
   U4315 : AO4 port map( A => n5129, B => n4413, C => n4738, D => n2134, Z => 
                           n2240);
   U4316 : AO7 port map( A => n5175, B => n5181, C => n4808, Z => n3616);
   U4317 : EON1 port map( A => n5049, B => n2577, C => n2646, D => n5230, Z => 
                           n2639);
   U4318 : AO2 port map( A => n5226, B => n2515, C => n5228, D => n2516, Z => 
                           n2513);
   U4319 : AO2 port map( A => n5217, B => n2922, C => n5224, D => n2924, Z => 
                           n2920);
   U4320 : AO4 port map( A => n2055, B => n4738, C => n5241, D => n4737, Z => 
                           n2286);
   U4321 : EO1 port map( A => n2147, B => n4769, C => n4738, D => n2147, Z => 
                           n2242);
   U4322 : AO2 port map( A => n5208, B => n3325, C => n5215, D => n3327, Z => 
                           n3323);
   U4323 : AO2 port map( A => n1888, B => n5199, C => n5197, D => n5140, Z => 
                           n2292);
   U4324 : AO2 port map( A => n5151, B => n5203, C => n5199, D => n2143, Z => 
                           n2138);
   U4325 : AO2 port map( A => n5198, B => n2015, C => n5240, D => n4507, Z => 
                           n2008);
   U4326 : AO2 port map( A => n2265, B => n5198, C => n5196, D => n1884, Z => 
                           n2347);
   U4327 : ND4 port map( A => n2307, B => n2308, C => n2309, D => n2310, Z => 
                           n1845);
   U4328 : AO2 port map( A => n5240, B => n5198, C => n5200, D => n2111, Z => 
                           n2308);
   U4329 : AO2 port map( A => n5203, B => n2311, C => n5202, D => n2312, Z => 
                           n2310);
   U4330 : AO2 port map( A => n5197, B => n2313, C => n2190, D => n5196, Z => 
                           n2309);
   U4331 : IVDA port map( A => n1762, Y => n_3417, Z => n4751);
   U4332 : IVDA port map( A => n1822, Y => n_3418, Z => n4747);
   U4333 : IVDA port map( A => n3295, Y => n_3419, Z => n4712);
   U4334 : AO2 port map( A => n2748, B => n4831, C => n2701, D => n5234, Z => 
                           n2747);
   U4335 : AO2 port map( A => n3155, B => n4815, C => n3108, D => n5223, Z => 
                           n3154);
   U4336 : AO2 port map( A => n3559, B => n4799, C => n3512, D => n5214, Z => 
                           n3558);
   U4337 : ND4 port map( A => n2136, B => n5122, C => n2138, D => n2139, Z => 
                           n2121);
   U4338 : AO2 port map( A => n2147, B => n5196, C => n2148, D => n5197, Z => 
                           n2136);
   U4339 : AO6 port map( A => n5201, B => n2140, C => n2141, Z => n2139);
   U4340 : IVI port map( A => n4356, Z => n4822);
   U4341 : IVI port map( A => n4808, Z => n4806);
   U4342 : IVI port map( A => n4839, Z => n4837);
   U4343 : IVI port map( A => n4356, Z => n4823);
   U4344 : IVI port map( A => n4808, Z => n4807);
   U4345 : AO2 port map( A => n5231, B => n5059, C => n4830, D => n2754, Z => 
                           n2792);
   U4346 : AO2 port map( A => n5220, B => n5237, C => n4814, D => n3161, Z => 
                           n3213);
   U4347 : AO2 port map( A => n5211, B => n5244, C => n4798, D => n3565, Z => 
                           n3617);
   U4348 : AO2 port map( A => n4770, B => n2225, C => n2110, D => n4515, Z => 
                           n2224);
   U4349 : AO2 port map( A => n5062, B => n5232, C => n5230, D => n2670, Z => 
                           n2851);
   U4350 : AO2 port map( A => n5103, B => n5221, C => n5219, D => n3078, Z => 
                           n3256);
   U4351 : AO2 port map( A => n5180, B => n5212, C => n5210, D => n3481, Z => 
                           n3661);
   U4352 : IVDA port map( A => n1762, Y => n_3420, Z => n4752);
   U4353 : IVDA port map( A => n1822, Y => n_3421, Z => n4748);
   U4354 : IVDA port map( A => n3295, Y => n_3422, Z => n4713);
   U4355 : IVI port map( A => n4381, Z => n4855);
   U4356 : IVI port map( A => n4381, Z => n4856);
   U4357 : IVI port map( A => n4839, Z => n4838);
   U4358 : EO1 port map( A => n2190, B => n4766, C => n4739, D => n2119, Z => 
                           n2228);
   U4359 : IVDA port map( A => n2060, Y => n4506, Z => n4736);
   U4360 : AO2 port map( A => n2749, B => n5231, C => n5046, D => n4839, Z => 
                           n2746);
   U4361 : AO2 port map( A => n3156, B => n5220, C => n5236, D => n4356, Z => 
                           n3153);
   U4362 : AO2 port map( A => n5127, B => n4515, C => n5137, D => n4767, Z => 
                           n2219);
   U4363 : AO2 port map( A => n3560, B => n5211, C => n5243, D => n4808, Z => 
                           n3557);
   U4364 : AO4 port map( A => n1001, B => n1002, C => n1003, D => n4927, Z => 
                           n1000);
   U4365 : AO4 port map( A => n1001, B => n4927, C => n1003, D => n1002, Z => 
                           n998);
   U4366 : AO4 port map( A => n191, B => n192_port, C => n193, D => n4946, Z =>
                           n190);
   U4367 : AO4 port map( A => n191, B => n4946, C => n193, D => n192_port, Z =>
                           n188);
   U4368 : AO4 port map( A => n4885, B => n270, C => n4368, D => n271, Z => 
                           n269);
   U4369 : AO4 port map( A => n4885, B => n1164, C => n4368, D => n1165, Z => 
                           n1163);
   U4370 : AO4 port map( A => n4885, B => n838, C => n4368, D => n839, Z => 
                           n837);
   U4371 : AO4 port map( A => n4885, B => n526, C => n4368, D => n527, Z => 
                           n525);
   U4372 : EON1 port map( A => n4368, B => n1221, C => n4370, D => n4668, Z => 
                           n1219);
   U4373 : ENI port map( A => n1237, B => n1238, Z => n4668);
   U4374 : AO4 port map( A => n4885, B => n932, C => n4368, D => n933, Z => 
                           n931);
   U4375 : AO4 port map( A => n4885, B => n113, C => n4368, D => n115, Z => 
                           n111);
   U4376 : AO4 port map( A => n4885, B => n1069, C => n4368, D => n1070, Z => 
                           n1068);
   U4377 : AO4 port map( A => n4885, B => n729, C => n4368, D => n730, Z => 
                           n728);
   U4378 : AO4 port map( A => n4885, B => n237, C => n4368, D => n238, Z => 
                           n236);
   U4379 : AO4 port map( A => n4885, B => n1042, C => n4368, D => n1043, Z => 
                           n1041);
   U4380 : AO4 port map( A => n4885, B => n700, C => n4368, D => n701, Z => 
                           n699);
   U4381 : AO4 port map( A => n4885, B => n398, C => n4368, D => n399, Z => 
                           n397);
   U4382 : AO4 port map( A => n4885, B => n208, C => n4368, D => n209, Z => 
                           n207);
   U4383 : AO4 port map( A => n4885, B => n1013, C => n4368, D => n1014, Z => 
                           n1012);
   U4384 : AO4 port map( A => n4885, B => n377, C => n4368, D => n378, Z => 
                           n376);
   U4385 : AO4 port map( A => n4885, B => n624, C => n4368, D => n625, Z => 
                           n623);
   U4386 : AO4 port map( A => n2195, B => n4737, C => n4736, D => n2196, Z => 
                           n2192);
   U4387 : AO3 port map( A => n5101, B => n2931, C => n2976, D => n2977, Z => 
                           n2974);
   U4388 : EO1 port map( A => n2989, B => n5225, C => n2991, D => n2936, Z => 
                           n2976);
   U4389 : AO4 port map( A => n2181, B => n2182, C => n4415, D => n2183, Z => 
                           n2176);
   U4390 : AO3 port map( A => n4736, B => n5141, C => n5132, D => n2187, Z => 
                           n2184);
   U4391 : IVDA port map( A => n3708, Y => n4352, Z => n4691);
   U4392 : AO7 port map( A => n4686, B => n4840, C => n4745, Z => n1938);
   U4393 : AO7 port map( A => n4687, B => n4840, C => n4746, Z => n1915);
   U4394 : AO7 port map( A => n4689, B => n4840, C => n4746, Z => n1908);
   U4395 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n4842, C => n4735, Z =>
                           n2459);
   U4396 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n4842, C => n4734, Z =>
                           n2455);
   U4397 : AO7 port map( A => n4669, B => n4842, C => n4735, Z => n2431);
   U4398 : AO7 port map( A => n4670, B => n4842, C => n4734, Z => n2427);
   U4399 : AO7 port map( A => n4671, B => n4842, C => n4735, Z => n2423);
   U4400 : AO3 port map( A => n5066, B => n4563, C => n2304, D => n2305, Z => 
                           n1507);
   U4401 : AO3 port map( A => n2078, B => n2057, C => n2314, D => n2315, Z => 
                           n2304);
   U4402 : AO2 port map( A => n5197, B => n2321, C => n1858, D => n5195, Z => 
                           n2314);
   U4403 : AO4 port map( A => n2076, B => n2077, C => n2050, D => n2078, Z => 
                           n2075);
   U4404 : AO2 port map( A => n2517, B => n4542, C => n2519, D => n2520, Z => 
                           n2512);
   U4405 : AO4 port map( A => n5098, B => n2984, C => n2985, D => n2986, Z => 
                           n2979);
   U4406 : AO2 port map( A => n2925, B => n4543, C => n2927, D => n2928, Z => 
                           n2919);
   U4407 : AO4 port map( A => n5155, B => n4738, C => n2290, D => n1882, Z => 
                           n2289);
   U4408 : AO6 port map( A => n2281, B => n4378, C => n4506, Z => n2290);
   U4409 : AO2 port map( A => n3328, B => n4544, C => n3330, D => n3331, Z => 
                           n3322);
   U4410 : AO7 port map( A => n3088, B => n3089, C => n5193, Z => n3080);
   U4411 : AO4 port map( A => n4823, B => n3090, C => n3091, D => n4715, Z => 
                           n3089);
   U4412 : AO4 port map( A => n5080, B => n3017, C => n4813, D => n3092, Z => 
                           n3088);
   U4413 : AO7 port map( A => n3491, B => n3492, C => n5206, Z => n3483);
   U4414 : AO4 port map( A => n4807, B => n3493, C => n3494, D => n4705, Z => 
                           n3492);
   U4415 : AO4 port map( A => n5157, B => n3420, C => n4797, D => n3495, Z => 
                           n3491);
   U4416 : AO3 port map( A => n5048, B => n2522, C => n2569, D => n2570, Z => 
                           n2568);
   U4417 : EO1 port map( A => n2583, B => n5229, C => n2585, D => n2526, Z => 
                           n2569);
   U4418 : AO4 port map( A => n2361, B => n4740, C => n2362, D => n1876, Z => 
                           n2360);
   U4419 : AO6 port map( A => n2146, B => n2196, C => n4737, Z => n2365);
   U4420 : AO4 port map( A => n2284, B => n1876, C => n2285, D => n4740, Z => 
                           n2283);
   U4421 : AO6 port map( A => n5150, B => n4769, C => n2289, Z => n2284);
   U4422 : AO3 port map( A => n5178, B => n3334, C => n3379, D => n3380, Z => 
                           n3377);
   U4423 : EO1 port map( A => n3392, B => n5216, C => n3394, D => n3339, Z => 
                           n3379);
   U4424 : IVDA port map( A => n1696, Y => n4543, Z => n4719);
   U4425 : IVDA port map( A => n2481, Y => n4544, Z => n4709);
   U4426 : AO3 port map( A => n5124, B => n4415, C => n2397, D => n2398, Z => 
                           n2395);
   U4427 : AO3 port map( A => n5241, B => n4412, C => n5070, D => n2405, Z => 
                           n2397);
   U4428 : AO2 port map( A => n5072, B => n2399, C => n4387, D => n2400, Z => 
                           n2398);
   U4429 : AO3 port map( A => n2323, B => n4740, C => n2324, D => n2325, Z => 
                           n2322);
   U4430 : ND3 port map( A => n2335, B => n5070, C => n2336, Z => n2324);
   U4431 : AO7 port map( A => n4685, B => n4850, C => n4733, Z => n2860);
   U4432 : AO7 port map( A => n4687, B => n4850, C => n4733, Z => n2782);
   U4433 : AO7 port map( A => n4680, B => n4850, C => n4723, Z => n3189);
   U4434 : AO7 port map( A => n4681, B => n4851, C => n4722, Z => n3145);
   U4435 : AO7 port map( A => n4678, B => n4844, C => n4758, Z => n1671);
   U4436 : AO7 port map( A => n4680, B => n4843, C => n4758, Z => n1641);
   U4437 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n4845, C => n4754, Z =>
                           n1757);
   U4438 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n4845, C => n4753, Z =>
                           n1753);
   U4439 : AO7 port map( A => n4669, B => n4844, C => n4754, Z => n1749);
   U4440 : AO7 port map( A => n4670, B => n4845, C => n4753, Z => n1745);
   U4441 : AO7 port map( A => n4671, B => n4845, C => n4754, Z => n1741);
   U4442 : ND4 port map( A => n2326, B => n2327, C => n2328, D => n2329, Z => 
                           n2325);
   U4443 : AO2 port map( A => n2332, B => n5151, C => n5154, D => n2334, Z => 
                           n2326);
   U4444 : EO1 port map( A => n2148, B => n5203, C => n2135, D => n2066, Z => 
                           n2328);
   U4445 : AO6 port map( A => n5072, B => n1873, C => n1874, Z => n1869);
   U4446 : AO4 port map( A => n1875, B => n1876, C => n4415, D => n1878, Z => 
                           n1874);
   U4447 : AO2 port map( A => n5235, B => n1887, C => n1888, D => n1881, Z => 
                           n1875);
   U4448 : AO7 port map( A => n2076, B => n2147, C => n2408, Z => n2407);
   U4449 : AO2 port map( A => n5198, B => n2134, C => n5142, D => n2409, Z => 
                           n2408);
   U4450 : AO7 port map( A => n2274, B => n5125, C => n2210, Z => n2409);
   U4451 : IVI port map( A => n2905, Z => n5220);
   U4452 : IVI port map( A => n3308, Z => n5211);
   U4453 : IVI port map( A => n3017, Z => n5223);
   U4454 : IVI port map( A => n3420, Z => n5214);
   U4455 : AO4 port map( A => n4736, B => n2068, C => n4739, D => n2367, Z => 
                           n2191);
   U4456 : AO6 port map( A => n2520, B => n2574, C => n4837, Z => n2770);
   U4457 : AO4 port map( A => n4727, B => n2585, C => n2593, D => n4827, Z => 
                           n2769);
   U4458 : AO6 port map( A => n2928, B => n2981, C => n4822, Z => n3177);
   U4459 : AO4 port map( A => n2905, B => n2991, C => n2999, D => n4812, Z => 
                           n3176);
   U4460 : AO6 port map( A => n3331, B => n3384, C => n4806, Z => n3581);
   U4461 : AO4 port map( A => n3308, B => n3394, C => n3402, D => n4796, Z => 
                           n3580);
   U4462 : AO4 port map( A => n2065, B => n2023, C => n5137, D => n2109, Z => 
                           n2350);
   U4463 : AO4 port map( A => n2119, B => n2066, C => n2076, D => n2241, Z => 
                           n2351);
   U4464 : AO4 port map( A => n2076, B => n2269, C => n2078, D => n2225, Z => 
                           n2267);
   U4465 : AO4 port map( A => n5153, B => n2116, C => n2263, D => n2066, Z => 
                           n2262);
   U4466 : EON1 port map( A => n2065, B => n2264, C => n5198, D => n2265, Z => 
                           n2261);
   U4467 : AO3 port map( A => n4413, B => n2216, C => n2278, D => n2279, Z => 
                           n2277);
   U4468 : IVI port map( A => n2109, Z => n5203);
   U4469 : ND4 port map( A => n2873, B => n2874, C => n2875, D => n2876, Z => 
                           n1958);
   U4470 : AO2 port map( A => n5230, B => n2610, C => n5226, D => n2544, Z => 
                           n2875);
   U4471 : AO2 port map( A => n4729, B => n5043, C => n5229, D => n5075, Z => 
                           n2873);
   U4472 : ND4 port map( A => n2810, B => n2811, C => n2812, D => n2813, Z => 
                           n1919);
   U4473 : AO2 port map( A => n5226, B => n2815, C => n5229, D => n2521, Z => 
                           n2811);
   U4474 : AO2 port map( A => n2701, B => n5232, C => n5230, D => n2614, Z => 
                           n2812);
   U4475 : AO2 port map( A => n5233, B => n5043, C => n5228, D => n2520, Z => 
                           n2810);
   U4476 : ND4 port map( A => n3285, B => n3286, C => n3287, D => n3288, Z => 
                           n1677);
   U4477 : AO2 port map( A => n5219, B => n3016, C => n5217, D => n2951, Z => 
                           n3287);
   U4478 : AO2 port map( A => n4716, B => n5095, C => n5225, D => n5100, Z => 
                           n3285);
   U4479 : ND4 port map( A => n3198, B => n3199, C => n3200, D => n3201, Z => 
                           n1648);
   U4480 : AO2 port map( A => n5217, B => n3204, C => n5225, D => n2930, Z => 
                           n3199);
   U4481 : AO2 port map( A => n3108, B => n5221, C => n5219, D => n3020, Z => 
                           n3200);
   U4482 : AO2 port map( A => n5222, B => n5095, C => n5224, D => n2928, Z => 
                           n3198);
   U4483 : ND4 port map( A => n3693, B => n3694, C => n3695, D => n3696, Z => 
                           n2462);
   U4484 : AO2 port map( A => n5210, B => n3419, C => n5208, D => n3354, Z => 
                           n3695);
   U4485 : AO2 port map( A => n4706, B => n5172, C => n5216, D => n5177, Z => 
                           n3693);
   U4486 : ND4 port map( A => n3602, B => n3603, C => n3604, D => n3605, Z => 
                           n2437);
   U4487 : AO2 port map( A => n5208, B => n3608, C => n5216, D => n3333, Z => 
                           n3603);
   U4488 : AO2 port map( A => n3512, B => n5212, C => n5210, D => n3423, Z => 
                           n3604);
   U4489 : AO2 port map( A => n5213, B => n5172, C => n5215, D => n3331, Z => 
                           n3602);
   U4490 : AO2 port map( A => n4770, B => n2188, C => n4766, D => n2189, Z => 
                           n2187);
   U4491 : EO1 port map( A => n2829, B => n2532, C => n2600, D => n4828, Z => 
                           n2828);
   U4492 : AO7 port map( A => n4397, B => n2684, C => n4837, Z => n2829);
   U4493 : EON1 port map( A => n1931, B => n4827, C => n1933, D => n5234, Z => 
                           n1927);
   U4494 : AO4 port map( A => n5053, B => n2577, C => n2578, D => n2579, Z => 
                           n2572);
   U4495 : EO1 port map( A => n3234, B => n1694, C => n3007, D => n4813, Z => 
                           n3233);
   U4496 : AO7 port map( A => n4395, B => n3092, C => n4822, Z => n3234);
   U4497 : EON1 port map( A => n1658, B => n4812, C => n2932, D => n5223, Z => 
                           n3193);
   U4498 : AO4 port map( A => n2985, B => n3049, C => n5115, D => n2931, Z => 
                           n3048);
   U4499 : EON1 port map( A => n2943, B => n3051, C => n4716, D => n3052, Z => 
                           n3047);
   U4500 : AO6 port map( A => n4813, B => n2998, C => n2999, Z => n2996);
   U4501 : AO4 port map( A => n2055, B => n4364, C => n4739, D => n2320, Z => 
                           n2364);
   U4502 : AO7 port map( A => n5139, B => n2076, C => n2116, Z => n2372);
   U4503 : EO1 port map( A => n3639, B => n2479, C => n3410, D => n4797, Z => 
                           n3638);
   U4504 : AO7 port map( A => n4371, B => n3495, C => n4806, Z => n3639);
   U4505 : EON1 port map( A => n2447, B => n4796, C => n3335, D => n5214, Z => 
                           n3597);
   U4506 : AO4 port map( A => n3388, B => n3452, C => n5192, D => n3334, Z => 
                           n3451);
   U4507 : EON1 port map( A => n3346, B => n3454, C => n4706, D => n3455, Z => 
                           n3450);
   U4508 : AO4 port map( A => n5175, B => n3387, C => n3388, D => n3389, Z => 
                           n3382);
   U4509 : AO2 port map( A => n5228, B => n2856, C => n2519, D => n2845, Z => 
                           n2852);
   U4510 : AO2 port map( A => n5204, B => n2789, C => n4400, D => n2790, Z => 
                           n2788);
   U4511 : AO3 port map( A => n2748, B => n4837, C => n2652, D => n2794, Z => 
                           n2789);
   U4512 : AO3 port map( A => n4725, B => n2646, C => n2791, D => n2792, Z => 
                           n2790);
   U4513 : AO2 port map( A => n4829, B => n2795, C => n5051, D => n5234, Z => 
                           n2794);
   U4514 : AO2 port map( A => n5224, B => n3261, C => n2927, D => n3250, Z => 
                           n3257);
   U4515 : AO2 port map( A => n5193, B => n3210, C => n4385, D => n3211, Z => 
                           n3209);
   U4516 : AO3 port map( A => n3155, B => n4822, C => n3060, D => n3214, Z => 
                           n3210);
   U4517 : AO3 port map( A => n4717, B => n3053, C => n3212, D => n3213, Z => 
                           n3211);
   U4518 : AO2 port map( A => n4814, B => n3215, C => n5090, D => n5223, Z => 
                           n3214);
   U4519 : AO4 port map( A => n2964, B => n4823, C => n5108, D => n4812, Z => 
                           n3093);
   U4520 : AO2 port map( A => n5217, B => n2960, C => n1658, D => n4716, Z => 
                           n2993);
   U4521 : AO2 port map( A => n5201, B => n2269, C => n5199, D => n2264, Z => 
                           n2307);
   U4522 : AO4 port map( A => n2210, B => n2032, C => n2273, D => n2274, Z => 
                           n2271);
   U4523 : AO2 port map( A => n5203, B => n2023, C => n5202, D => n5153, Z => 
                           n2006);
   U4524 : AO2 port map( A => n2018, B => n5200, C => n5201, D => n2021, Z => 
                           n2007);
   U4525 : AO2 port map( A => n5215, B => n3666, C => n3330, D => n3655, Z => 
                           n3662);
   U4526 : AO2 port map( A => n5206, B => n3614, C => n4386, D => n3615, Z => 
                           n3613);
   U4527 : AO3 port map( A => n3559, B => n4806, C => n3463, D => n3618, Z => 
                           n3614);
   U4528 : AO3 port map( A => n4707, B => n3456, C => n3616, D => n3617, Z => 
                           n3615);
   U4529 : AO2 port map( A => n4798, B => n3619, C => n5167, D => n5214, Z => 
                           n3618);
   U4530 : AO4 port map( A => n3367, B => n4807, C => n5185, D => n4796, Z => 
                           n3496);
   U4531 : AO4 port map( A => n5037, B => n4731, C => n1961, D => n4730, Z => 
                           n1959);
   U4532 : AO6 port map( A => n1954, B => n1962, C => n1963, Z => n1961);
   U4533 : AO4 port map( A => n4838, B => n1964, C => n5049, D => n4727, Z => 
                           n1963);
   U4534 : AO2 port map( A => n4521, B => n2826, C => n4400, D => n2827, Z => 
                           n2825);
   U4535 : AO3 port map( A => n4725, B => n2532, C => n2830, D => n5039, Z => 
                           n2826);
   U4536 : AO7 port map( A => n4728, B => n2731, C => n2828, Z => n2827);
   U4537 : AO4 port map( A => n2840, B => n4730, C => n2841, D => n4731, Z => 
                           n2839);
   U4538 : AO6 port map( A => n2521, B => n2708, C => n4837, Z => n2847);
   U4539 : AO2 port map( A => n4521, B => n2744, C => n4400, D => n2745, Z => 
                           n2743);
   U4540 : AO3 port map( A => n4827, B => n2532, C => n2750, D => n2751, Z => 
                           n2744);
   U4541 : AO3 port map( A => n2755, B => n2522, C => n2756, D => n2757, Z => 
                           n2741);
   U4542 : AO2 port map( A => n2760, B => n5230, C => n4729, D => n2761, Z => 
                           n2756);
   U4543 : AO2 port map( A => n5228, B => n2758, C => n5052, D => n2519, Z => 
                           n2757);
   U4544 : AO3 port map( A => n1933, B => n2522, C => n2771, D => n2772, Z => 
                           n2762);
   U4545 : AO2 port map( A => n5229, B => n2778, C => n5041, D => n4729, Z => 
                           n2771);
   U4546 : AO4 port map( A => n2493, B => n4731, C => n2494, D => n4730, Z => 
                           n2492);
   U4547 : AO6 port map( A => n2495, B => n4397, C => n2497, Z => n2494);
   U4548 : AO6 port map( A => n4833, B => n2501, C => n2502, Z => n2493);
   U4549 : AO4 port map( A => n5058, B => n4728, C => n2499, D => n4838, Z => 
                           n2497);
   U4550 : AO4 port map( A => n5086, B => n4720, C => n3278, D => n4721, Z => 
                           n3277);
   U4551 : AO6 port map( A => n1684, B => n1682, C => n3279, Z => n3278);
   U4552 : AO4 port map( A => n4822, B => n1685, C => n5080, D => n4715, Z => 
                           n3279);
   U4553 : AO2 port map( A => n4520, B => n3231, C => n4385, D => n3232, Z => 
                           n3230);
   U4554 : AO3 port map( A => n4717, B => n1694, C => n3235, D => n5094, Z => 
                           n3231);
   U4555 : AO7 port map( A => n4714, B => n3137, C => n3233, Z => n3232);
   U4556 : AO4 port map( A => n3245, B => n4721, C => n3246, D => n4720, Z => 
                           n3244);
   U4557 : AO6 port map( A => n2930, B => n3114, C => n4822, Z => n3252);
   U4558 : AO2 port map( A => n4520, B => n3151, C => n4385, D => n3152, Z => 
                           n3150);
   U4559 : AO3 port map( A => n4812, B => n1694, C => n3157, D => n3158, Z => 
                           n3151);
   U4560 : AO3 port map( A => n3162, B => n2931, C => n3163, D => n3164, Z => 
                           n3148);
   U4561 : AO2 port map( A => n3167, B => n5219, C => n4716, D => n3168, Z => 
                           n3163);
   U4562 : AO2 port map( A => n5224, B => n3165, C => n5091, D => n2927, Z => 
                           n3164);
   U4563 : AO3 port map( A => n2932, B => n2931, C => n3178, D => n3179, Z => 
                           n3169);
   U4564 : AO2 port map( A => n5225, B => n3185, C => n5102, D => n4716, Z => 
                           n3178);
   U4565 : AO4 port map( A => n2898, B => n4720, C => n2900, D => n4721, Z => 
                           n2897);
   U4566 : AO6 port map( A => n2902, B => n4395, C => n2903, Z => n2900);
   U4567 : AO6 port map( A => n4818, B => n2908, C => n2909, Z => n2898);
   U4568 : AO4 port map( A => n5096, B => n4714, C => n2906, D => n4822, Z => 
                           n2903);
   U4569 : AO2 port map( A => n1888, B => n2355, C => n5120, D => n5198, Z => 
                           n2353);
   U4570 : AO7 port map( A => n2196, B => n2274, C => n2210, Z => n2355);
   U4571 : AO2 port map( A => n5072, B => n2217, C => n5070, D => n2218, Z => 
                           n2207);
   U4572 : AO3 port map( A => n4377, B => n2222, C => n2223, D => n2224, Z => 
                           n2217);
   U4573 : AO2 port map( A => n5149, B => n4770, C => n2165, D => n4765, Z => 
                           n2220);
   U4574 : AO4 port map( A => n2042, B => n1876, C => n2043, D => n4740, Z => 
                           n2041);
   U4575 : AO6 port map( A => n4767, B => n2046, C => n2047, Z => n2043);
   U4576 : AO4 port map( A => n4378, B => n5125, C => n2059, D => n4736, Z => 
                           n2053);
   U4577 : AO4 port map( A => n5163, B => n4710, C => n3686, D => n4711, Z => 
                           n3685);
   U4578 : AO6 port map( A => n2469, B => n2467, C => n3687, Z => n3686);
   U4579 : AO4 port map( A => n4806, B => n2470, C => n5157, D => n4705, Z => 
                           n3687);
   U4580 : AO2 port map( A => n4522, B => n3636, C => n4386, D => n3637, Z => 
                           n3635);
   U4581 : AO3 port map( A => n4707, B => n2479, C => n3640, D => n5171, Z => 
                           n3636);
   U4582 : AO7 port map( A => n4704, B => n3541, C => n3638, Z => n3637);
   U4583 : AO4 port map( A => n3650, B => n4711, C => n3651, D => n4710, Z => 
                           n3649);
   U4584 : AO6 port map( A => n3333, B => n3518, C => n4806, Z => n3657);
   U4585 : AO2 port map( A => n4522, B => n3555, C => n4386, D => n3556, Z => 
                           n3554);
   U4586 : AO3 port map( A => n4796, B => n2479, C => n3561, D => n3562, Z => 
                           n3555);
   U4587 : AO3 port map( A => n3566, B => n3334, C => n3567, D => n3568, Z => 
                           n3552);
   U4588 : AO2 port map( A => n3571, B => n5210, C => n4706, D => n3572, Z => 
                           n3567);
   U4589 : AO2 port map( A => n5215, B => n3569, C => n5168, D => n3330, Z => 
                           n3568);
   U4590 : AO3 port map( A => n3335, B => n3334, C => n3582, D => n3583, Z => 
                           n3573);
   U4591 : AO2 port map( A => n5216, B => n3589, C => n5179, D => n4706, Z => 
                           n3582);
   U4592 : AO4 port map( A => n3301, B => n4710, C => n3303, D => n4711, Z => 
                           n3300);
   U4593 : AO6 port map( A => n3305, B => n4371, C => n3306, Z => n3303);
   U4594 : AO6 port map( A => n4802, B => n3311, C => n3312, Z => n3301);
   U4595 : AO4 port map( A => n5173, B => n4704, C => n3309, D => n4806, Z => 
                           n3306);
   U4596 : AO4 port map( A => n5138, B => n1843, C => n1844, D => n1845, Z => 
                           n1841);
   U4597 : AO3 port map( A => n5131, B => n4519, C => n1848, D => n5071, Z => 
                           n1843);
   U4598 : IVDA port map( A => n1949, Y => n4542, Z => n4724);
   U4599 : AO3 port map( A => n4728, B => n2612, C => n2867, D => n2868, Z => 
                           n2866);
   U4600 : AO7 port map( A => n2869, B => n4839, C => n5048, Z => n2868);
   U4601 : AO3 port map( A => n2905, B => n3018, C => n3282, D => n3283, Z => 
                           n3281);
   U4602 : AO7 port map( A => n3284, B => n4356, C => n5101, Z => n3283);
   U4603 : AO3 port map( A => n4739, B => n2225, C => n2317, D => n2318, Z => 
                           n2316);
   U4604 : AO2 port map( A => n2319, B => n4504, C => n4507, D => n2072, Z => 
                           n2318);
   U4605 : AO3 port map( A => n3308, B => n3421, C => n3690, D => n3691, Z => 
                           n3689);
   U4606 : AO7 port map( A => n3692, B => n4808, C => n5178, Z => n3691);
   U4607 : AO3 port map( A => n2786, B => n2536, C => n2787, D => n2788, Z => 
                           n2785);
   U4608 : AO7 port map( A => n2797, B => n2798, C => n4521, Z => n2787);
   U4609 : AO3 port map( A => n3207, B => n2945, C => n3208, D => n3209, Z => 
                           n3206);
   U4610 : AO7 port map( A => n3218, B => n3219, C => n4520, Z => n3208);
   U4611 : AO3 port map( A => n3611, B => n3348, C => n3612, D => n3613, Z => 
                           n3610);
   U4612 : AO7 port map( A => n3622, B => n3623, C => n4522, Z => n3612);
   U4613 : AO4 port map( A => n4726, B => n2642, C => n5045, D => n4827, Z => 
                           n2842);
   U4614 : AO4 port map( A => n4718, B => n3049, C => n5115, D => n4812, Z => 
                           n3247);
   U4615 : AO4 port map( A => n2145, B => n2066, C => n2065, D => n2034, Z => 
                           n2144);
   U4616 : AO4 port map( A => n2055, B => n4739, C => n4737, D => n2057, Z => 
                           n2054);
   U4617 : AO4 port map( A => n4708, B => n3452, C => n5192, D => n4796, Z => 
                           n3652);
   U4618 : ND4 port map( A => n2292, B => n2293, C => n2294, D => n2295, Z => 
                           n2282);
   U4619 : AO2 port map( A => n2296, B => n5200, C => n5203, D => n2297, Z => 
                           n2295);
   U4620 : AO2 port map( A => n5201, B => n2189, C => n5127, D => n5202, Z => 
                           n2294);
   U4621 : AO2 port map( A => n5198, B => n5119, C => n5134, D => n5196, Z => 
                           n2293);
   U4622 : AO2 port map( A => n2134, B => n4515, C => n4767, D => n2071, Z => 
                           n2403);
   U4623 : AO2 port map( A => n4504, B => n5119, C => n4766, D => n5140, Z => 
                           n2404);
   U4624 : EO1 port map( A => n5143, B => n4507, C => n2199, D => n4737, Z => 
                           n2198);
   U4625 : AO2 port map( A => n4769, B => n2200, C => n4767, D => n1884, Z => 
                           n2197);
   U4626 : AO4 port map( A => n2679, B => n1966, C => n2495, D => n4837, Z => 
                           n2832);
   U4627 : AO4 port map( A => n3087, B => n4715, C => n2902, D => n4822, Z => 
                           n3237);
   U4628 : AO4 port map( A => n3490, B => n4705, C => n3305, D => n4806, Z => 
                           n3642);
   U4629 : AO6 port map( A => n3083, B => n3084, C => n2945, Z => n3082);
   U4630 : AO2 port map( A => n5223, B => n5102, C => n3087, D => n4816, Z => 
                           n3083);
   U4631 : AO2 port map( A => n3049, B => n4356, C => n3085, D => n5220, Z => 
                           n3084);
   U4632 : AO4 port map( A => n2109, B => n2110, C => n2111, D => n2070, Z => 
                           n2108);
   U4633 : AO6 port map( A => n3486, B => n3487, C => n3348, Z => n3485);
   U4634 : AO2 port map( A => n5214, B => n5179, C => n3490, D => n4800, Z => 
                           n3486);
   U4635 : AO2 port map( A => n3452, B => n4808, C => n3488, D => n5211, Z => 
                           n3487);
   U4636 : ND3 port map( A => n1657, B => n4395, C => n1696, Z => n2988);
   U4637 : IVI port map( A => n1966, Z => n5231);
   U4638 : IVI port map( A => n2611, Z => n5234);
   U4639 : AO4 port map( A => n5035, B => n4837, C => n5046, D => n1966, Z => 
                           n2766);
   U4640 : AO4 port map( A => n5106, B => n4822, C => n5236, D => n4715, Z => 
                           n3173);
   U4641 : AO4 port map( A => n5183, B => n4806, C => n5243, D => n4705, Z => 
                           n3577);
   U4642 : AO4 port map( A => n4728, B => n2553, C => n4828, D => n2628, Z => 
                           n2626);
   U4643 : NR3 port map( A => n4838, B => n5074, C => n5063, Z => n2627);
   U4644 : AO4 port map( A => n4714, B => n2961, C => n4813, D => n3035, Z => 
                           n3033);
   U4645 : NR3 port map( A => n4823, B => n5097, C => n5088, Z => n3034);
   U4646 : AO4 port map( A => n4704, B => n3364, C => n4797, D => n3438, Z => 
                           n3436);
   U4647 : NR3 port map( A => n4807, B => n5174, C => n5165, Z => n3437);
   U4648 : IVDA port map( A => n1473, Y => n4545, Z => n4694);
   U4649 : NR4 port map( A => n1464, B => n4695, C => n4693, D => n4696, Z => 
                           n1463);
   U4650 : ND4 port map( A => n4545, B => n4699, C => n4698, D => n4428, Z => 
                           n1464);
   U4651 : AO4 port map( A => n2848, B => n4827, C => n2611, D => n2849, Z => 
                           n2846);
   U4652 : AO4 port map( A => n3253, B => n4812, C => n3017, D => n3254, Z => 
                           n3251);
   U4653 : AO4 port map( A => n3658, B => n4796, C => n3420, D => n3659, Z => 
                           n3656);
   U4654 : AO4 port map( A => n2068, B => n4412, C => n2133, D => n4736, Z => 
                           n2239);
   U4655 : AO2 port map( A => n2583, B => n5231, C => n4839, D => n2582, Z => 
                           n2751);
   U4656 : AO2 port map( A => n2679, B => n4397, C => n5076, D => n4360, Z => 
                           n2712);
   U4657 : AO6 port map( A => n4828, B => n2592, C => n2593, Z => n2590);
   U4658 : AO2 port map( A => n2989, B => n5220, C => n4356, D => n1657, Z => 
                           n3158);
   U4659 : AO2 port map( A => n3087, B => n4395, C => n5087, D => n4355, Z => 
                           n3118);
   U4660 : EON1 port map( A => n4412, B => n2021, C => n4765, D => n2018, Z => 
                           n2339);
   U4661 : AO4 port map( A => n1857, B => n2142, C => n4378, D => n2130, Z => 
                           n2141);
   U4662 : AO2 port map( A => n3392, B => n5211, C => n4808, D => n2446, Z => 
                           n3562);
   U4663 : AO2 port map( A => n3490, B => n4371, C => n5164, D => n4358, Z => 
                           n3522);
   U4664 : AO6 port map( A => n4797, B => n3401, C => n3402, Z => n3399);
   U4665 : AO2 port map( A => n5061, B => n5233, C => n5230, D => n2801, Z => 
                           n2886);
   U4666 : AO7 port map( A => n2680, B => n2681, C => n5204, Z => n2672);
   U4667 : AO4 port map( A => n4838, B => n2682, C => n2683, D => n1966, Z => 
                           n2681);
   U4668 : AO4 port map( A => n5049, B => n2611, C => n4828, D => n2684, Z => 
                           n2680);
   U4669 : AO4 port map( A => n2556, B => n4838, C => n5077, D => n4827, Z => 
                           n2685);
   U4670 : AO2 port map( A => n5226, B => n2552, C => n1931, D => n4729, Z => 
                           n2587);
   U4671 : AO2 port map( A => n5105, B => n5222, C => n5219, D => n3222, Z => 
                           n3271);
   U4672 : AO4 port map( A => n4412, B => n2164, C => n4737, D => n2168, Z => 
                           n2167);
   U4673 : AO2 port map( A => n5182, B => n5213, C => n5210, D => n3626, Z => 
                           n3679);
   U4674 : AO2 port map( A => n5208, B => n3363, C => n2447, D => n4706, Z => 
                           n3396);
   U4675 : AO7 port map( A => n2698, B => n2699, C => n5205, Z => n2697);
   U4676 : AO4 port map( A => n4725, B => n2600, C => n4827, D => n2702, Z => 
                           n2698);
   U4677 : AO4 port map( A => n4838, B => n2700, C => n2701, D => n4727, Z => 
                           n2699);
   U4678 : AO7 port map( A => n5031, B => n2549, C => n5234, Z => n2547);
   U4679 : AO4 port map( A => n5064, B => n4731, C => n4730, D => n2550, Z => 
                           n2549);
   U4680 : AO2 port map( A => n2501, B => n5204, C => n2552, D => n5205, Z => 
                           n2551);
   U4681 : AO7 port map( A => n2530, B => n2531, C => n4839, Z => n2529);
   U4682 : AO4 port map( A => n2533, B => n2534, C => n5056, D => n2536, Z => 
                           n2530);
   U4683 : AO4 port map( A => n4731, B => n2532, C => n4542, D => n4730, Z => 
                           n2531);
   U4684 : AO7 port map( A => n3105, B => n3106, C => n5194, Z => n3104);
   U4685 : AO4 port map( A => n4717, B => n3007, C => n4813, D => n3109, Z => 
                           n3105);
   U4686 : AO4 port map( A => n4823, B => n3107, C => n3108, D => n2905, Z => 
                           n3106);
   U4687 : AO7 port map( A => n5082, B => n2957, C => n5223, Z => n2955);
   U4688 : AO4 port map( A => n5089, B => n4720, C => n4721, D => n2958, Z => 
                           n2957);
   U4689 : AO2 port map( A => n2908, B => n5193, C => n2960, D => n5194, Z => 
                           n2959);
   U4690 : AO7 port map( A => n2940, B => n2941, C => n4356, Z => n2939);
   U4691 : AO4 port map( A => n2942, B => n2943, C => n5239, D => n2945, Z => 
                           n2940);
   U4692 : AO4 port map( A => n4720, B => n1694, C => n4543, D => n4721, Z => 
                           n2941);
   U4693 : AO6 port map( A => n2131, B => n2132, C => n4740, Z => n2122);
   U4694 : AO2 port map( A => n4515, B => n2021, C => n4767, D => n2135, Z => 
                           n2131);
   U4695 : AO2 port map( A => n4770, B => n2133, C => n2134, D => n4765, Z => 
                           n2132);
   U4696 : AO7 port map( A => n3509, B => n3510, C => n5207, Z => n3508);
   U4697 : AO4 port map( A => n4707, B => n3410, C => n4797, D => n3513, Z => 
                           n3509);
   U4698 : AO4 port map( A => n4807, B => n3511, C => n3512, D => n3308, Z => 
                           n3510);
   U4699 : AO7 port map( A => n5159, B => n3360, C => n5214, Z => n3358);
   U4700 : AO4 port map( A => n5166, B => n4710, C => n4711, D => n3361, Z => 
                           n3360);
   U4701 : AO2 port map( A => n3311, B => n5206, C => n3363, D => n5207, Z => 
                           n3362);
   U4702 : AO7 port map( A => n3343, B => n3344, C => n4808, Z => n3342);
   U4703 : AO4 port map( A => n3345, B => n3346, C => n5246, D => n3348, Z => 
                           n3343);
   U4704 : AO4 port map( A => n4710, B => n2479, C => n4544, D => n4711, Z => 
                           n3344);
   U4705 : IVDA port map( A => n2102, Y => n4507, Z => n4738);
   U4706 : AO4 port map( A => n2735, B => n2611, C => n4837, D => n2649, Z => 
                           n2799);
   U4707 : AO4 port map( A => n3141, B => n3017, C => n4822, D => n3057, Z => 
                           n3220);
   U4708 : AO4 port map( A => n3545, B => n3420, C => n4806, D => n3460, Z => 
                           n3624);
   U4709 : AO3 port map( A => n5083, B => n4813, C => n4385, D => n3072, Z => 
                           n3070);
   U4710 : AO6 port map( A => n3065, B => n3076, C => n4718, Z => n3075);
   U4711 : AO3 port map( A => n5160, B => n4797, C => n4386, D => n3475, Z => 
                           n3473);
   U4712 : AO6 port map( A => n3468, B => n3479, C => n4708, Z => n3478);
   U4713 : AO7 port map( A => n4686, B => n4855, C => n4751, Z => n1783);
   U4714 : AO7 port map( A => n4687, B => n4855, C => n4752, Z => n1779);
   U4715 : AO7 port map( A => n4689, B => n4855, C => n4752, Z => n1772);
   U4716 : AO7 port map( A => n4678, B => n4856, C => n4750, Z => n1817);
   U4717 : AO7 port map( A => n4680, B => n4855, C => n4750, Z => n1809);
   U4718 : AO7 port map( A => n4681, B => n4855, C => n4749, Z => n1804);
   U4719 : AO7 port map( A => n4673, B => n4856, C => n4748, Z => n1866);
   U4720 : AO7 port map( A => n4674, B => n4856, C => n4748, Z => n1839);
   U4721 : AO6 port map( A => n2675, B => n2676, C => n2536, Z => n2674);
   U4722 : AO2 port map( A => n5234, B => n5041, C => n2679, D => n4832, Z => 
                           n2675);
   U4723 : AO2 port map( A => n2642, B => n4839, C => n2677, D => n5231, Z => 
                           n2676);
   U4724 : ND3 port map( A => n2582, B => n4397, C => n1949, Z => n2581);
   U4725 : ND3 port map( A => n2446, B => n4371, C => n2481, Z => n3391);
   U4726 : IVDA port map( A => n1924, Y => n4400, Z => n4731);
   U4727 : IVDA port map( A => n2899, Y => n4385, Z => n4720);
   U4728 : IVDA port map( A => n3302, Y => n4386, Z => n4710);
   U4729 : IVDA port map( A => n1466, Y => n_3423, Z => n4693);
   U4730 : IVDA port map( A => n1467, Y => n_3424, Z => n4696);
   U4731 : IVDA port map( A => n1477, Y => n_3425, Z => n4700);
   U4732 : IVDA port map( A => n2049, Y => n4504, Z => n4737);
   U4733 : IVDA port map( A => n2056, Y => n4515, Z => n4739);
   U4734 : AO4 port map( A => n2582, B => n4726, C => n4827, D => n2731, Z => 
                           n2797);
   U4735 : AO4 port map( A => n4837, B => n2525, C => n2645, D => n4728, Z => 
                           n2798);
   U4736 : EON1 port map( A => n2534, B => n2644, C => n4729, D => n2645, Z => 
                           n2640);
   U4737 : AO4 port map( A => n2578, B => n2642, C => n5045, D => n2522, Z => 
                           n2641);
   U4738 : AO4 port map( A => n1657, B => n4718, C => n4812, D => n3137, Z => 
                           n3218);
   U4739 : AO4 port map( A => n4822, B => n2935, C => n3052, D => n4715, Z => 
                           n3219);
   U4740 : EO1 port map( A => n5151, B => n4404, C => n2200, D => n4737, Z => 
                           n2335);
   U4741 : AO4 port map( A => n2446, B => n4708, C => n4796, D => n3541, Z => 
                           n3622);
   U4742 : AO4 port map( A => n4806, B => n3338, C => n3455, D => n4705, Z => 
                           n3623);
   U4743 : AO2 port map( A => n2854, B => n4729, C => n5226, D => n2855, Z => 
                           n2853);
   U4744 : EO1 port map( A => n5229, B => n2544, C => n2815, D => n2522, Z => 
                           n2850);
   U4745 : AO2 port map( A => n3259, B => n4716, C => n5217, D => n3260, Z => 
                           n3258);
   U4746 : EO1 port map( A => n5225, B => n2951, C => n3204, D => n2931, Z => 
                           n3255);
   U4747 : AO2 port map( A => n5144, B => n4768, C => n5143, D => n4504, Z => 
                           n2227);
   U4748 : AO7 port map( A => n4378, B => n2093, C => n5070, Z => n2166);
   U4749 : AO2 port map( A => n3664, B => n4706, C => n5208, D => n3665, Z => 
                           n3663);
   U4750 : EO1 port map( A => n5216, B => n3354, C => n3608, D => n3334, Z => 
                           n3660);
   U4751 : AO3 port map( A => n4837, B => n2642, C => n4400, D => n2733, Z => 
                           n2715);
   U4752 : AO6 port map( A => n5035, B => n5231, C => n2734, Z => n2733);
   U4753 : AO4 port map( A => n4827, B => n2574, C => n2735, D => n2611, Z => 
                           n2734);
   U4754 : AO6 port map( A => n2556, B => n4400, C => n2558, Z => n2545);
   U4755 : AO4 port map( A => n4730, B => n2559, C => n5044, D => n2533, Z => 
                           n2558);
   U4756 : AO3 port map( A => n4822, B => n3049, C => n4385, D => n3139, Z => 
                           n3121);
   U4757 : AO6 port map( A => n5106, B => n5220, C => n3140, Z => n3139);
   U4758 : AO4 port map( A => n4812, B => n2981, C => n3141, D => n3017, Z => 
                           n3140);
   U4759 : AO6 port map( A => n2964, B => n4385, C => n2965, Z => n2952);
   U4760 : AO4 port map( A => n4721, B => n2966, C => n5104, D => n2942, Z => 
                           n2965);
   U4761 : AO3 port map( A => n4806, B => n3452, C => n4386, D => n3543, Z => 
                           n3525);
   U4762 : AO6 port map( A => n5183, B => n5211, C => n3544, Z => n3543);
   U4763 : AO4 port map( A => n4796, B => n3384, C => n3545, D => n3420, Z => 
                           n3544);
   U4764 : AO6 port map( A => n3367, B => n4386, C => n3368, Z => n3355);
   U4765 : AO4 port map( A => n4711, B => n3369, C => n5181, D => n3345, Z => 
                           n3368);
   U4766 : AO6 port map( A => n4387, B => n1892, C => n4563, Z => n1868);
   U4767 : AO2 port map( A => n2445, B => n2446, C => n2447, D => n4802, Z => 
                           n2444);
   U4768 : AO2 port map( A => n1926, B => n2582, C => n1931, D => n4829, Z => 
                           n2805);
   U4769 : AO2 port map( A => n1656, B => n1657, C => n1658, D => n4818, Z => 
                           n1655);
   U4770 : AO4 port map( A => n5035, B => n4837, C => n2749, D => n4727, Z => 
                           n2843);
   U4771 : EON1 port map( A => n2647, B => n1966, C => n2801, D => n4834, Z => 
                           n2800);
   U4772 : AO4 port map( A => n5106, B => n4822, C => n3156, D => n2905, Z => 
                           n3248);
   U4773 : EON1 port map( A => n3055, B => n2905, C => n3222, D => n4820, Z => 
                           n3221);
   U4774 : AO4 port map( A => n5183, B => n4806, C => n3560, D => n3308, Z => 
                           n3653);
   U4775 : EON1 port map( A => n3458, B => n3308, C => n3626, D => n4804, Z => 
                           n3625);
   U4776 : AO4 port map( A => n2611, B => n2721, C => n4827, D => n1964, Z => 
                           n2720);
   U4777 : AO4 port map( A => n3017, B => n3127, C => n4812, D => n1685, Z => 
                           n3126);
   U4778 : AO4 port map( A => n3420, B => n3531, C => n4796, D => n2470, Z => 
                           n3530);
   U4779 : IVDA port map( A => n3708, Y => n4353, Z => n4692);
   U4780 : AO3 port map( A => n5050, B => n4828, C => n4400, D => n2664, Z => 
                           n2662);
   U4781 : AO6 port map( A => n2657, B => n2668, C => n4726, Z => n2667);
   U4782 : IVDA port map( A => n2044, Y => n4387, Z => n4740);
   U4783 : ND3 port map( A => n5036, B => n4360, C => n5205, Z => n2546);
   U4784 : ND3 port map( A => n5111, B => n4355, C => n5194, Z => n2954);
   U4785 : ND3 port map( A => n5188, B => n4357, C => n5207, Z => n3357);
   U4786 : IVI port map( A => n4394, Z => n4858);
   U4787 : IVI port map( A => n4889, Z => n4886);
   U4788 : AO2 port map( A => n1330, B => n1331, C => n4916, D => n1332, Z => 
                           n1278);
   U4789 : AO2 port map( A => n4911, B => n998, C => n999, D => n1000, Z => 
                           n970);
   U4790 : AO2 port map( A => n4957, B => n188, C => n189, D => n190, Z => n145
                           );
   U4791 : AO3 port map( A => n4888, B => n4484, C => n299, D => n300, Z => 
                           n4047);
   U4792 : AO6 port map( A => n301, B => n4790, C => n302, Z => n300);
   U4793 : AO2 port map( A => n4784, B => n323, C => n324, D => n4787, Z => 
                           n299);
   U4794 : AO4 port map( A => n4885, B => n303, C => n4368, D => n304, Z => 
                           n302);
   U4795 : AO3 port map( A => n4887, B => n4485, C => n754, D => n755, Z => 
                           n4053);
   U4796 : AO6 port map( A => n756, B => n4789, C => n757, Z => n755);
   U4797 : AO2 port map( A => n4783, B => n782, C => n783, D => n4788, Z => 
                           n754);
   U4798 : AO4 port map( A => n4885, B => n758, C => n4368, D => n759, Z => 
                           n757);
   U4799 : AO3 port map( A => n4886, B => n4486, C => n1101, D => n1102, Z => 
                           n4059);
   U4800 : AO6 port map( A => n1103, B => n4789, C => n1104, Z => n1102);
   U4801 : AO2 port map( A => n4783, B => n1145, C => n1146, D => n4788, Z => 
                           n1101);
   U4802 : AO4 port map( A => n4885, B => n1105, C => n4368, D => n1106, Z => 
                           n1104);
   U4803 : AO3 port map( A => n4887, B => n4487, C => n497, D => n498, Z => 
                           n4065);
   U4804 : AO6 port map( A => n499, B => n4790, C => n500, Z => n498);
   U4805 : AO2 port map( A => n4784, B => n515, C => n516, D => n4787, Z => 
                           n497);
   U4806 : AO4 port map( A => n4885, B => n501, C => n4368, D => n502, Z => 
                           n500);
   U4807 : AO4 port map( A => n4885, B => n468, C => n4368, D => n469, Z => 
                           n467);
   U4808 : AO3 port map( A => n4887, B => n4482, C => n594, D => n595, Z => 
                           n4034);
   U4809 : AO6 port map( A => n596, B => n4790, C => n597, Z => n595);
   U4810 : AO2 port map( A => n4784, B => n613, C => n614, D => n4787, Z => 
                           n594);
   U4811 : AO3 port map( A => n4887, B => n4483, C => n792, D => n793, Z => 
                           n4041);
   U4812 : AO6 port map( A => n794, B => n4789, C => n795, Z => n793);
   U4813 : AO2 port map( A => n4783, B => n822, C => n823, D => n4788, Z => 
                           n792);
   U4814 : ND3 port map( A => n4886, B => n5010, C => n1301, Z => n163);
   U4815 : ND3 port map( A => n1315, B => n4886, C => n5021, Z => n164);
   U4816 : IVDA port map( A => v_KEY_COLUMN_21_port, Y => n4576, Z => n4682);
   U4817 : IVDA port map( A => v_KEY_COLUMN_22_port, Y => n4577, Z => n4683);
   U4818 : IVDA port map( A => v_KEY_COLUMN_13_port, Y => n4392, Z => n4676);
   U4819 : AO4 port map( A => n4885, B => n565, C => n4368, D => n566, Z => 
                           n564);
   U4820 : AO4 port map( A => n4885, B => n598, C => n4368, D => n599, Z => 
                           n597);
   U4821 : AO4 port map( A => n4885, B => n796, C => n4368, D => n797, Z => 
                           n795);
   U4822 : AO4 port map( A => n4885, B => n891, C => n4368, D => n892, Z => 
                           n890);
   U4823 : AO4 port map( A => n4885, B => n427, C => n4368, D => n428, Z => 
                           n426);
   U4824 : AO3 port map( A => n4886, B => n4479, C => n1216, D => n1217, Z => 
                           n4016);
   U4825 : AO6 port map( A => n1218, B => n4789, C => n1219, Z => n1217);
   U4826 : AO2 port map( A => n4783, B => n1263, C => n1264, D => n4788, Z => 
                           n1216);
   U4827 : IVDA port map( A => v_KEY_COLUMN_16_port, Y => n4454, Z => n4678);
   U4828 : IVDA port map( A => v_KEY_COLUMN_10_port, Y => n4569, Z => n4674);
   U4829 : IVDA port map( A => v_KEY_COLUMN_30_port, Y => n4567, Z => n4690);
   U4830 : IVDA port map( A => v_KEY_COLUMN_18_port, Y => n4456, Z => n4680);
   U4831 : IVDA port map( A => v_KEY_COLUMN_23_port, Y => n4458, Z => n4684);
   U4832 : IVDA port map( A => v_KEY_COLUMN_14_port, Y => n4571, Z => n4677);
   U4833 : IVDA port map( A => v_KEY_COLUMN_8_port, Y => n4391, Z => n4673);
   U4834 : AO4 port map( A => n1302, B => n163, C => n164, D => n1303, Z => 
                           n1281);
   U4835 : AO4 port map( A => n982, B => n163, C => n164, D => n983, Z => n973)
                           ;
   U4836 : AO4 port map( A => n162, B => n163, C => n164, D => n165, Z => n149)
                           ;
   U4837 : AO7 port map( A => n5011, B => n4471, C => n1436, Z => n1434);
   U4838 : AO4 port map( A => v_RAM_OUT0_9_port, B => n2153, C => n2154, D => 
                           n4563, Z => n1492);
   U4839 : IVDA port map( A => v_KEY_COLUMN_24_port, Y => n4565, Z => n4685);
   U4840 : AO6 port map( A => n3058, B => n3059, C => n4403, Z => n3043);
   U4841 : NR4 port map( A => n3045, B => n3046, C => n3047, D => n3048, Z => 
                           n3044);
   U4842 : AO2 port map( A => v_RAM_OUT0_17_port, B => n3063, C => n5110, D => 
                           n5222, Z => n3058);
   U4843 : AO6 port map( A => n3461, B => n3462, C => n4401, Z => n3446);
   U4844 : NR4 port map( A => n3448, B => n3449, C => n3450, D => n3451, Z => 
                           n3447);
   U4845 : AO2 port map( A => v_RAM_OUT0_1_port, B => n3466, C => n5187, D => 
                           n5213, Z => n3461);
   U4846 : IVDA port map( A => v_KEY_COLUMN_26_port, Y => n4389, Z => n4687);
   U4847 : IVDA port map( A => v_KEY_COLUMN_27_port, Y => n4566, Z => n4688);
   U4848 : IVDA port map( A => v_KEY_COLUMN_17_port, Y => n4455, Z => n4679);
   U4849 : IVDA port map( A => v_KEY_COLUMN_19_port, Y => n4457, Z => n4681);
   U4850 : IVDA port map( A => v_KEY_COLUMN_2_port, Y => n4459, Z => n4669);
   U4851 : IVDA port map( A => v_KEY_COLUMN_3_port, Y => n4460, Z => n4670);
   U4852 : IVDA port map( A => v_KEY_COLUMN_7_port, Y => n4568, Z => n4672);
   U4853 : IVDA port map( A => v_KEY_COLUMN_25_port, Y => n4375, Z => n4686);
   U4854 : AO4 port map( A => n2970, B => n2971, C => n2972, D => n4564, Z => 
                           n1618);
   U4855 : AO3 port map( A => n3026, B => n2945, C => n3027, D => n4564, Z => 
                           n2970);
   U4856 : AO2 port map( A => n4782, B => n2973, C => n2974, D => n4402, Z => 
                           n2972);
   U4857 : AO4 port map( A => n3040, B => n3041, C => v_RAM_OUT0_23_port, D => 
                           n3042, Z => n3039);
   U4858 : AO3 port map( A => n3079, B => n4721, C => n3080, D => n5081, Z => 
                           n3040);
   U4859 : AO4 port map( A => n3443, B => n3444, C => v_RAM_OUT0_7_port, D => 
                           n3445, Z => n3442);
   U4860 : AO3 port map( A => n3482, B => n4711, C => n3483, D => n5158, Z => 
                           n3443);
   U4861 : AO3 port map( A => n1606, B => n1893, C => n1939, D => n1940, Z => 
                           n4035);
   U4862 : AO7 port map( A => n4685, B => n4840, C => n4746, Z => n1941);
   U4863 : AO3 port map( A => n1590, B => n1893, C => n1909, D => n1910, Z => 
                           n4134);
   U4864 : AO7 port map( A => n4688, B => n4840, C => n4745, Z => n1911);
   U4865 : AO3 port map( A => n5033, B => n1893, C => n1902, D => n1903, Z => 
                           n4166);
   U4866 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n4840, C => n4745, Z 
                           => n1904);
   U4867 : AO3 port map( A => n1575, B => n1893, C => n1899, D => n1900, Z => 
                           n4167);
   U4868 : AO7 port map( A => n4690, B => n4840, C => n4746, Z => n1901);
   U4869 : AO3 port map( A => n1568, B => n1893, C => n1894, D => n1895, Z => 
                           n4168);
   U4870 : AO7 port map( A => v_KEY_COLUMN_31_port, B => n4840, C => n4745, Z 
                           => n1897);
   U4871 : AO3 port map( A => n1813, B => n1967, C => n1993, D => n1994, Z => 
                           n4169);
   U4872 : AO7 port map( A => n4678, B => n4841, C => n4744, Z => n1995);
   U4873 : AO3 port map( A => n1663, B => n1967, C => n1989, D => n1990, Z => 
                           n4170);
   U4874 : AO7 port map( A => n4679, B => n4841, C => n4743, Z => n1992);
   U4875 : AO3 port map( A => n1805, B => n1967, C => n1985, D => n1986, Z => 
                           n4171);
   U4876 : AO7 port map( A => n4680, B => n4841, C => n4744, Z => n1988);
   U4877 : AO3 port map( A => n1632, B => n1967, C => n1981, D => n1982, Z => 
                           n4172);
   U4878 : AO7 port map( A => n4681, B => n4840, C => n4743, Z => n1984);
   U4879 : AO3 port map( A => n1628, B => n1967, C => n1978, D => n1979, Z => 
                           n4173);
   U4880 : AO7 port map( A => v_KEY_COLUMN_20_port, B => n4840, C => n4744, Z 
                           => n1980);
   U4881 : AO3 port map( A => n1611, B => n1967, C => n1968, D => n1969, Z => 
                           n4176);
   U4882 : AO7 port map( A => n4684, B => n4840, C => n4743, Z => n1971);
   U4883 : AO3 port map( A => n1517, B => n1997, C => n2373, D => n2374, Z => 
                           n4177);
   U4884 : AO7 port map( A => n4673, B => n4840, C => n4742, Z => n2375);
   U4885 : AO3 port map( A => n1512, B => n1997, C => n2340, D => n2341, Z => 
                           n4178);
   U4886 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n4841, C => n4741, Z =>
                           n2342);
   U4887 : AO3 port map( A => n1507, B => n1997, C => n2301, D => n2302, Z => 
                           n4179);
   U4888 : AO7 port map( A => n4674, B => n4841, C => n4742, Z => n2303);
   U4889 : AO3 port map( A => n1502, B => n1997, C => n2252, D => n2253, Z => 
                           n4180);
   U4890 : AO7 port map( A => n4675, B => n4841, C => n4741, Z => n2254);
   U4891 : AO3 port map( A => n1498, B => n1997, C => n2201, D => n2202, Z => 
                           n4181);
   U4892 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n4841, C => n4742, Z 
                           => n2203);
   U4893 : AO3 port map( A => n1492, B => n1997, C => n2149, D => n2150, Z => 
                           n4182);
   U4894 : AO7 port map( A => n4676, B => n4841, C => n4741, Z => n2152);
   U4895 : AO3 port map( A => n1487, B => n1997, C => n2079, D => n2080, Z => 
                           n4183);
   U4896 : AO7 port map( A => n4677, B => n4841, C => n4742, Z => n2081);
   U4897 : AO3 port map( A => n1480, B => n1997, C => n1998, D => n1999, Z => 
                           n4184);
   U4898 : AO7 port map( A => v_KEY_COLUMN_15_port, B => n4841, C => n4741, Z 
                           => n2000);
   U4899 : AO3 port map( A => n2456, B => n2410, C => n2457, D => n2458, Z => 
                           n4185);
   U4900 : AO2 port map( A => n2460, B => n4580, C => v_RAM_OUT0_7_port, D => 
                           n2461, Z => n2456);
   U4901 : AO3 port map( A => n2428, B => n2410, C => n2429, D => n2430, Z => 
                           n4187);
   U4902 : AO2 port map( A => v_RAM_OUT0_7_port, B => n2433, C => n5161, D => 
                           n4580, Z => n2428);
   U4903 : AO3 port map( A => n1531, B => n2410, C => n2415, D => n2416, Z => 
                           n4191);
   U4904 : AO7 port map( A => v_KEY_COLUMN_6_port, B => n4841, C => n4735, Z =>
                           n2417);
   U4905 : AO3 port map( A => n1524, B => n2410, C => n2411, D => n2412, Z => 
                           n4192);
   U4906 : AO7 port map( A => n4672, B => n4842, C => n4734, Z => n2413);
   U4907 : AO3 port map( A => n2857, B => n2483, C => n2858, D => n2859, Z => 
                           n4193);
   U4908 : AO2 port map( A => n2862, B => n4579, C => v_RAM_OUT0_31_port, D => 
                           n2863, Z => n2857);
   U4909 : AO3 port map( A => n1601, B => n2483, C => n2817, D => n2818, Z => 
                           n4194);
   U4910 : AO7 port map( A => n4686, B => n4850, C => n4732, Z => n2820);
   U4911 : AO3 port map( A => n2779, B => n2483, C => n2780, D => n2781, Z => 
                           n4195);
   U4912 : AO2 port map( A => v_RAM_OUT0_31_port, B => n2784, C => n5030, D => 
                           n4579, Z => n2779);
   U4913 : AO3 port map( A => n1590, B => n2483, C => n2736, D => n2737, Z => 
                           n4196);
   U4914 : AO7 port map( A => n4688, B => n4850, C => n4732, Z => n2738);
   U4915 : AO3 port map( A => n1584, B => n2483, C => n2689, D => n2690, Z => 
                           n4197);
   U4916 : AO7 port map( A => n4689, B => n4850, C => n4733, Z => n2692);
   U4917 : AO3 port map( A => n5033, B => n2483, C => n2629, D => n2630, Z => 
                           n4198);
   U4918 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n4850, C => n4732, Z 
                           => n2631);
   U4919 : AO3 port map( A => n1575, B => n2483, C => n2561, D => n2562, Z => 
                           n4199);
   U4920 : AO7 port map( A => n4690, B => n4850, C => n4733, Z => n2563);
   U4921 : AO3 port map( A => n1568, B => n2483, C => n2484, D => n2485, Z => 
                           n4200);
   U4922 : AO7 port map( A => v_KEY_COLUMN_31_port, B => n4850, C => n4732, Z 
                           => n2486);
   U4923 : AO3 port map( A => n1813, B => n2888, C => n3262, D => n3263, Z => 
                           n4201);
   U4924 : AO7 port map( A => n4678, B => n4851, C => n4723, Z => n3264);
   U4925 : AO3 port map( A => n1663, B => n2888, C => n3223, D => n3224, Z => 
                           n4202);
   U4926 : AO7 port map( A => n4679, B => n4851, C => n4722, Z => n3225);
   U4927 : AO3 port map( A => n1628, B => n2888, C => n3097, D => n3098, Z => 
                           n4205);
   U4928 : AO7 port map( A => v_KEY_COLUMN_20_port, B => n4851, C => n4723, Z 
                           => n3099);
   U4929 : AO3 port map( A => n5065, B => n2888, C => n3036, D => n3037, Z => 
                           n4206);
   U4930 : AO7 port map( A => n4682, B => n4850, C => n4722, Z => n3038);
   U4931 : AO3 port map( A => n1618, B => n2888, C => n2967, D => n2968, Z => 
                           n4207);
   U4932 : AO7 port map( A => n4683, B => n4850, C => n4723, Z => n2969);
   U4933 : AO3 port map( A => n1611, B => n2888, C => n2889, D => n2890, Z => 
                           n4208);
   U4934 : AO7 port map( A => n4684, B => n4850, C => n4722, Z => n2891);
   U4935 : AO3 port map( A => n1481, B => n1492, C => n1493, D => n1494, Z => 
                           n4214);
   U4936 : AO7 port map( A => n4676, B => n4849, C => n1486, Z => n1497);
   U4937 : AO3 port map( A => n1525, B => n1562, C => n1563, D => n1564, Z => 
                           n4217);
   U4938 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n4850, C => n4760, Z =>
                           n1566);
   U4939 : AO3 port map( A => n1525, B => n1557, C => n1558, D => n1559, Z => 
                           n4218);
   U4940 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n4850, C => n4759, Z =>
                           n1561);
   U4941 : AO3 port map( A => n1525, B => n1551, C => n1552, D => n1553, Z => 
                           n4219);
   U4942 : AO7 port map( A => n4669, B => n4849, C => n4760, Z => n1556);
   U4943 : AO3 port map( A => n1525, B => n1545, C => n1546, D => n1547, Z => 
                           n4220);
   U4944 : AO7 port map( A => n4670, B => n4849, C => n4759, Z => n1550);
   U4945 : AO3 port map( A => n1525, B => n1539, C => n1540, D => n1541, Z => 
                           n4221);
   U4946 : AO7 port map( A => n4671, B => n4849, C => n4760, Z => n1544);
   U4947 : AO3 port map( A => n5073, B => n1525, C => n1536, D => n1537, Z => 
                           n4222);
   U4948 : AO7 port map( A => v_KEY_COLUMN_5_port, B => n4849, C => n4759, Z =>
                           n1538);
   U4949 : AO3 port map( A => n1525, B => n1531, C => n1532, D => n1533, Z => 
                           n4223);
   U4950 : AO7 port map( A => v_KEY_COLUMN_6_port, B => n4849, C => n4760, Z =>
                           n1534);
   U4951 : AO3 port map( A => n1524, B => n1525, C => n1526, D => n1527, Z => 
                           n4224);
   U4952 : AO7 port map( A => n4672, B => n4849, C => n4759, Z => n1529);
   U4953 : AO3 port map( A => n1492, B => n1698, C => n1706, D => n1707, Z => 
                           n4246);
   U4954 : AO7 port map( A => n4676, B => n4844, C => n4755, Z => n1709);
   U4955 : AO3 port map( A => n1492, B => n1818, C => n1826, D => n1827, Z => 
                           n4278);
   U4956 : AO7 port map( A => n4676, B => n4856, C => n4747, Z => n1829);
   U4957 : EON1 port map( A => n4633, B => n1435, C => n4633, D => n1434, Z => 
                           n4290);
   U4958 : AO4 port map( A => n2488, B => n2489, C => v_RAM_OUT0_31_port, D => 
                           n2490, Z => n1568);
   U4959 : AO3 port map( A => n2528, B => n4728, C => n2529, D => 
                           v_RAM_OUT0_31_port, Z => n2489);
   U4960 : AO3 port map( A => n2545, B => n4828, C => n2546, D => n2547, Z => 
                           n2488);
   U4961 : AO6 port map( A => v_RAM_OUT0_29_port, B => n2491, C => n2492, Z => 
                           n2490);
   U4962 : AO4 port map( A => n2893, B => n2894, C => v_RAM_OUT0_23_port, D => 
                           n2895, Z => n1611);
   U4963 : AO3 port map( A => n2938, B => n4714, C => n2939, D => 
                           v_RAM_OUT0_23_port, Z => n2894);
   U4964 : AO3 port map( A => n2952, B => n4812, C => n2954, D => n2955, Z => 
                           n2893);
   U4965 : AO6 port map( A => n4782, B => n2896, C => n2897, Z => n2895);
   U4966 : AO3 port map( A => n2343, B => n4563, C => n2344, D => n2345, Z => 
                           n1512);
   U4967 : ND4 port map( A => n5067, B => n2346, C => n2347, D => n2348, Z => 
                           n2345);
   U4968 : ND4 port map( A => n5071, B => n2352, C => n2353, D => n2354, Z => 
                           n2344);
   U4969 : AO6 port map( A => v_RAM_OUT0_15_port, B => n2359, C => n2360, Z => 
                           n2343);
   U4970 : AO7 port map( A => n2255, B => n4563, C => n2256, Z => n1502);
   U4971 : AO2 port map( A => n2257, B => n2258, C => n2259, D => n2260, Z => 
                           n2256);
   U4972 : AO6 port map( A => v_RAM_OUT0_15_port, B => n2282, C => n2283, Z => 
                           n2255);
   U4973 : AO4 port map( A => n3296, B => n3297, C => v_RAM_OUT0_7_port, D => 
                           n3298, Z => n1524);
   U4974 : AO3 port map( A => n3341, B => n4704, C => n3342, D => 
                           v_RAM_OUT0_7_port, Z => n3297);
   U4975 : AO3 port map( A => n3355, B => n4796, C => n3357, D => n3358, Z => 
                           n3296);
   U4976 : AO6 port map( A => v_RAM_OUT0_5_port, B => n3299, C => n3300, Z => 
                           n3298);
   U4977 : AO4 port map( A => n2033, B => n2076, C => n2065, D => n1889, Z => 
                           n2330);
   U4978 : AO7 port map( A => v_RAM_OUT0_9_port, B => n2082, C => n2083_port, Z
                           => n1487);
   U4979 : AO3 port map( A => n2084_port, B => n2085_port, C => 
                           v_RAM_OUT0_9_port, D => n2086_port, Z => n2083_port)
                           ;
   U4980 : AO3 port map( A => n2078, B => n5142, C => v_RAM_OUT0_15_port, D => 
                           n5121, Z => n2085_port);
   U4981 : IVDA port map( A => v_KEY_COLUMN_28_port, Y => n4390, Z => n4689);
   U4982 : IVDA port map( A => v_KEY_COLUMN_11_port, Y => n4570, Z => n4675);
   U4983 : IVDA port map( A => v_KEY_COLUMN_4_port, Y => n4461, Z => n4671);
   U4984 : AO4 port map( A => n2525, B => n2526, C => v_RAM_OUT0_25_port, D => 
                           n5042, Z => n2507);
   U4985 : AO4 port map( A => n2521, B => n2522, C => n1933, D => n4516, Z => 
                           n2508);
   U4986 : AO3 port map( A => n5035, B => n2511, C => n2512, D => n2513, Z => 
                           n2509);
   U4987 : AO4 port map( A => n2935, B => n2936, C => v_RAM_OUT0_17_port, D => 
                           n5085, Z => n2914);
   U4988 : AO4 port map( A => n2930, B => n2931, C => n2932, D => n4517, Z => 
                           n2915);
   U4989 : AO3 port map( A => n5106, B => n2918, C => n2919, D => n2920, Z => 
                           n2916);
   U4990 : AO4 port map( A => n3338, B => n3339, C => v_RAM_OUT0_1_port, D => 
                           n5162, Z => n3317);
   U4991 : AO4 port map( A => n3333, B => n3334, C => n3335, D => n4518, Z => 
                           n3318);
   U4992 : AO3 port map( A => n5183, B => n3321, C => n3322, D => n3323, Z => 
                           n3319);
   U4993 : AO4 port map( A => n4395, B => n3065, C => v_RAM_OUT0_18_port, D => 
                           n3066, Z => n3063);
   U4994 : AO2 port map( A => n3067, B => n1696, C => n5103, D => n4780, Z => 
                           n3066);
   U4995 : AO4 port map( A => n4371, B => n3468, C => v_RAM_OUT0_2_port, D => 
                           n3469, Z => n3466);
   U4996 : AO2 port map( A => n3470, B => n2481, C => n5180, D => n4779, Z => 
                           n3469);
   U4997 : AO3 port map( A => n1697, B => n4823, C => n3060, D => n3061, Z => 
                           n3059);
   U4998 : AO4 port map( A => n4378, B => n1889, C => v_RAM_OUT0_10_port, D => 
                           n1890, Z => n1887);
   U4999 : AO3 port map( A => n2482, B => n4807, C => n3463, D => n3464, Z => 
                           n3462);
   U5000 : AO6 port map( A => n2124, B => n2125, C => n1876, Z => n2123);
   U5001 : AO2 port map( A => n4770, B => n2127, C => n4507, D => n2128, Z => 
                           n2125);
   U5002 : EO1 port map( A => n1890, B => n4769, C => n2130, D => n4365, Z => 
                           n2124);
   U5003 : AO3 port map( A => n2112, B => n2065, C => n2113, D => n2114, Z => 
                           n2084_port);
   U5004 : AO2 port map( A => n2117, B => n5126, C => n2119, D => n5199, Z => 
                           n2113);
   U5005 : EO1 port map( A => n5145, B => n5197, C => n2077, D => n2116, Z => 
                           n2114);
   U5006 : AO7 port map( A => v_RAM_OUT0_9_port, B => n5068, C => n2378, Z => 
                           n1517);
   U5007 : AO3 port map( A => n2182, B => n1873, C => n2379, D => n2380, Z => 
                           n2378);
   U5008 : AO6 port map( A => n5128, B => n4387, C => n4563, Z => n2380);
   U5009 : AO2 port map( A => n5070, B => n2385, C => v_RAM_OUT0_15_port, D => 
                           n2386, Z => n2379);
   U5010 : AO4 port map( A => n2564, B => n2565, C => n2566, D => n4579, Z => 
                           n1575);
   U5011 : AO3 port map( A => n2619, B => n2536, C => n2620, D => n4579, Z => 
                           n2564);
   U5012 : AO2 port map( A => v_RAM_OUT0_29_port, B => n2567, C => n2568, D => 
                           n4379, Z => n2566);
   U5013 : AO4 port map( A => v_RAM_OUT0_9_port, B => n2002, C => n2003, D => 
                           n4563, Z => n1480);
   U5014 : AO2 port map( A => v_RAM_OUT0_15_port, B => n2004, C => n2005, D => 
                           n4415, Z => n2003);
   U5015 : AO6 port map( A => n2039, B => n2040, C => n2041, Z => n2002);
   U5016 : ND4 port map( A => n2006, B => n2007, C => n2008, D => n2009, Z => 
                           n2005);
   U5017 : AO4 port map( A => n3373, B => n3374, C => n3375, D => n4580, Z => 
                           n1531);
   U5018 : AO3 port map( A => n3429, B => n3348, C => n3430, D => n4580, Z => 
                           n3373);
   U5019 : AO2 port map( A => v_RAM_OUT0_5_port, B => n3376, C => n3377, D => 
                           n4401, Z => n3375);
   U5020 : EON1 port map( A => n1880, B => n1881, C => n1882, D => n1881, Z => 
                           n1879);
   U5021 : AO2 port map( A => n5137, B => v_RAM_OUT0_10_port, C => n1884, D => 
                           n4378, Z => n1880);
   U5022 : AO3 port map( A => n1481, B => n1517, C => n1518, D => n1519, Z => 
                           n4209);
   U5023 : AO7 port map( A => n4673, B => n4849, C => n1486, Z => n1522);
   U5024 : AO3 port map( A => n1481, B => n1512, C => n1513, D => n1514, Z => 
                           n4210);
   U5025 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n4849, C => n1486, Z =>
                           n1516);
   U5026 : AO3 port map( A => n1481, B => n1507, C => n1508, D => n1509, Z => 
                           n4211);
   U5027 : AO7 port map( A => n4674, B => n4849, C => n1486, Z => n1511);
   U5028 : AO3 port map( A => n1481, B => n1502, C => n1503, D => n1504, Z => 
                           n4212);
   U5029 : AO7 port map( A => n4675, B => n4849, C => n1486, Z => n1506);
   U5030 : AO3 port map( A => n1481, B => n1498, C => n1499, D => n1500, Z => 
                           n4213);
   U5031 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n4849, C => n1486, Z 
                           => n1501);
   U5032 : AO3 port map( A => n1481, B => n1487, C => n1488, D => n1489, Z => 
                           n4215);
   U5033 : AO7 port map( A => n4677, B => n4849, C => n1486, Z => n1491);
   U5034 : AO3 port map( A => n1480, B => n1481, C => n1482, D => n1483, Z => 
                           n4216);
   U5035 : AO7 port map( A => v_KEY_COLUMN_15_port, B => n4849, C => n1486, Z 
                           => n1485);
   U5036 : AO3 port map( A => n1569, B => n1606, C => n1607, D => n1608, Z => 
                           n4225);
   U5037 : AO7 port map( A => n4685, B => n4843, C => n1574, Z => n1610);
   U5038 : AO3 port map( A => n1569, B => n1601, C => n1602, D => n1603, Z => 
                           n4226);
   U5039 : AO7 port map( A => n4686, B => n4843, C => n1574, Z => n1605);
   U5040 : AO3 port map( A => n1569, B => n1595, C => n1596, D => n1597, Z => 
                           n4227);
   U5041 : AO7 port map( A => n4687, B => n4843, C => n1574, Z => n1600);
   U5042 : AO3 port map( A => n1569, B => n1590, C => n1591, D => n1592, Z => 
                           n4228);
   U5043 : AO7 port map( A => n4688, B => n4843, C => n1574, Z => n1594);
   U5044 : AO3 port map( A => n1569, B => n1584, C => n1585, D => n1586, Z => 
                           n4229);
   U5045 : AO7 port map( A => n4689, B => n4843, C => n1574, Z => n1589);
   U5046 : AO3 port map( A => n5033, B => n1569, C => n1581, D => n1582, Z => 
                           n4230);
   U5047 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n4843, C => n1574, Z 
                           => n1583);
   U5048 : AO3 port map( A => n1569, B => n1575, C => n1576, D => n1577, Z => 
                           n4231);
   U5049 : AO7 port map( A => n4690, B => n4843, C => n1574, Z => n1579);
   U5050 : AO3 port map( A => n1568, B => n1569, C => n1570, D => n1571, Z => 
                           n4232);
   U5051 : AO7 port map( A => v_KEY_COLUMN_31_port, B => n4843, C => n1574, Z 
                           => n1573);
   U5052 : AO3 port map( A => n1668, B => n1612, C => n1669, D => n1670, Z => 
                           n4233);
   U5053 : AO2 port map( A => n1675, B => n4564, C => v_RAM_OUT0_23_port, D => 
                           n1676, Z => n1668);
   U5054 : AO3 port map( A => n1612, B => n1663, C => n1664, D => n1665, Z => 
                           n4234);
   U5055 : AO7 port map( A => n4679, B => n4844, C => n4757, Z => n1667);
   U5056 : AO3 port map( A => n1638, B => n1612, C => n1639, D => n1640, Z => 
                           n4235);
   U5057 : AO2 port map( A => v_RAM_OUT0_23_port, B => n1644, C => n5084, D => 
                           n4564, Z => n1638);
   U5058 : AO3 port map( A => n1612, B => n1632, C => n1633, D => n1634, Z => 
                           n4236);
   U5059 : AO7 port map( A => n4681, B => n4843, C => n4757, Z => n1637);
   U5060 : AO3 port map( A => n1612, B => n1628, C => n1629, D => n1630, Z => 
                           n4237);
   U5061 : AO7 port map( A => v_KEY_COLUMN_20_port, B => n4843, C => n4758, Z 
                           => n1631);
   U5062 : AO3 port map( A => n5065, B => n1612, C => n1624, D => n1625, Z => 
                           n4238);
   U5063 : AO7 port map( A => n4682, B => n4843, C => n4757, Z => n1627);
   U5064 : AO3 port map( A => n1612, B => n1618, C => n1619, D => n1620, Z => 
                           n4239);
   U5065 : AO7 port map( A => n4683, B => n4843, C => n4758, Z => n1622);
   U5066 : AO3 port map( A => n1611, B => n1612, C => n1613, D => n1614, Z => 
                           n4240);
   U5067 : AO7 port map( A => n4684, B => n4843, C => n4757, Z => n1616);
   U5068 : AO3 port map( A => n1517, B => n1698, C => n1722, D => n1723, Z => 
                           n4241);
   U5069 : AO7 port map( A => n4673, B => n4844, C => n4756, Z => n1725);
   U5070 : AO3 port map( A => n1512, B => n1698, C => n1719, D => n1720, Z => 
                           n4242);
   U5071 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n4844, C => n4755, Z =>
                           n1721);
   U5072 : AO3 port map( A => n1507, B => n1698, C => n1716, D => n1717, Z => 
                           n4243);
   U5073 : AO7 port map( A => n4674, B => n4844, C => n4756, Z => n1718);
   U5074 : AO3 port map( A => n1502, B => n1698, C => n1713, D => n1714, Z => 
                           n4244);
   U5075 : AO7 port map( A => n4675, B => n4844, C => n4755, Z => n1715);
   U5076 : AO3 port map( A => n1498, B => n1698, C => n1710, D => n1711, Z => 
                           n4245);
   U5077 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n4844, C => n4756, Z 
                           => n1712);
   U5078 : AO3 port map( A => n1487, B => n1698, C => n1703, D => n1704, Z => 
                           n4247);
   U5079 : AO7 port map( A => n4677, B => n4844, C => n4756, Z => n1705);
   U5080 : AO3 port map( A => n1480, B => n1698, C => n1699, D => n1700, Z => 
                           n4248);
   U5081 : AO7 port map( A => v_KEY_COLUMN_15_port, B => n4844, C => n4755, Z 
                           => n1701);
   U5082 : AO3 port map( A => n5073, B => n1727, C => n1735, D => n1736, Z => 
                           n4254);
   U5083 : AO7 port map( A => v_KEY_COLUMN_5_port, B => n4844, C => n4753, Z =>
                           n1737);
   U5084 : AO3 port map( A => n1531, B => n1727, C => n1732, D => n1733, Z => 
                           n4255);
   U5085 : AO7 port map( A => v_KEY_COLUMN_6_port, B => n4844, C => n4754, Z =>
                           n1734);
   U5086 : AO3 port map( A => n1524, B => n1727, C => n1728, D => n1729, Z => 
                           n4256);
   U5087 : AO7 port map( A => n4672, B => n4844, C => n4753, Z => n1730);
   U5088 : AO3 port map( A => n1575, B => n1758, C => n1763, D => n1764, Z => 
                           n4263);
   U5089 : AO7 port map( A => n4690, B => n4855, C => n4752, Z => n1765);
   U5090 : AO3 port map( A => n1568, B => n1758, C => n1759, D => n1760, Z => 
                           n4264);
   U5091 : AO7 port map( A => v_KEY_COLUMN_31_port, B => n4855, C => n4751, Z 
                           => n1761);
   U5092 : AO3 port map( A => n1618, B => n1787, C => n1792, D => n1793, Z => 
                           n4271);
   U5093 : AO7 port map( A => n4683, B => n4855, C => n4750, Z => n1794);
   U5094 : AO3 port map( A => n1611, B => n1787, C => n1788, D => n1789, Z => 
                           n4272);
   U5095 : AO7 port map( A => n4684, B => n4855, C => n4749, Z => n1790);
   U5096 : AO3 port map( A => n1863, B => n1818, C => n1864, D => n1865, Z => 
                           n4273);
   U5097 : AO2 port map( A => n1868, B => n1869, C => n5068, D => n4563, Z => 
                           n1863);
   U5098 : AO3 port map( A => n1512, B => n1818, C => n1859, D => n1860, Z => 
                           n4274);
   U5099 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n4856, C => n4747, Z =>
                           n1862);
   U5100 : AO3 port map( A => n1502, B => n1818, C => n1833, D => n1834, Z => 
                           n4276);
   U5101 : AO7 port map( A => n4675, B => n4856, C => n4747, Z => n1835);
   U5102 : AO3 port map( A => n1487, B => n1818, C => n1823, D => n1824, Z => 
                           n4279);
   U5103 : AO7 port map( A => n4677, B => n4856, C => n4748, Z => n1825);
   U5104 : AO3 port map( A => n1480, B => n1818, C => n1819, D => n1820, Z => 
                           n4280);
   U5105 : AO7 port map( A => v_KEY_COLUMN_15_port, B => n4856, C => n4747, Z 
                           => n1821);
   U5106 : AO3 port map( A => n1531, B => n3291, C => n3370, D => n3371, Z => 
                           n4287);
   U5107 : AO7 port map( A => v_KEY_COLUMN_6_port, B => n4856, C => n4713, Z =>
                           n3372);
   U5108 : AO3 port map( A => n1524, B => n3291, C => n3292, D => n3293, Z => 
                           n4288);
   U5109 : AO7 port map( A => n4672, B => n4856, C => n4712, Z => n3294);
   U5110 : ND4 port map( A => n2368, B => n2369, C => n2370, D => n2371, Z => 
                           n2359);
   U5111 : AO2 port map( A => n5203, B => n2145, C => n5130, D => n5202, Z => 
                           n2370);
   U5112 : AO2 port map( A => n2372, B => n2033, C => n5143, D => n5200, Z => 
                           n2371);
   U5113 : ND4 port map( A => n2169, B => n2170, C => n2171, D => n2172, Z => 
                           n2155);
   U5114 : AO2 port map( A => n5151, B => n5198, C => n5200, D => n2173, Z => 
                           n2172);
   U5115 : AO2 port map( A => n5202, B => n5135, C => n2147, D => n5196, Z => 
                           n2170);
   U5116 : AO2 port map( A => n5199, B => n2069, C => n5197, D => n2077, Z => 
                           n2169);
   U5117 : ND4 port map( A => n2026, B => n2027, C => n2028, D => n2029, Z => 
                           n2004);
   U5118 : AO2 port map( A => n5200, B => n2033, C => n5203, D => n2034, Z => 
                           n2028);
   U5119 : AO2 port map( A => n2030, B => n5242, C => n5202, D => n2032, Z => 
                           n2029);
   U5120 : AO2 port map( A => n5198, B => n1889, C => n5196, D => n2035, Z => 
                           n2027);
   U5121 : NR3 port map( A => n1418, B => n5009, C => n5011, Z => n1409);
   U5122 : ND4 port map( A => v_RAM_OUT0_9_port, B => n2206, C => n2207, D => 
                           n2208, Z => n2205);
   U5123 : AO3 port map( A => n2233, B => n4415, C => n2234, D => n2235, Z => 
                           n2204);
   U5124 : ND4 port map( A => n2227, B => n4387, C => n2228, D => n2229, Z => 
                           n2206);
   U5125 : IVI port map( A => n4889, Z => n4887);
   U5126 : AO2 port map( A => v_RAM_OUT0_12_port, B => n5140, C => n4404, D => 
                           n2145, Z => n1858);
   U5127 : AO3 port map( A => n4737, B => n2241, C => n2231, D => n2242, Z => 
                           n2236);
   U5128 : AO7 port map( A => n2239, B => n2240, C => n5070, Z => n2238);
   U5129 : IVDA port map( A => n2524, Y => n4516, Z => n4729);
   U5130 : IVDA port map( A => n2934, Y => n4517, Z => n4716);
   U5131 : IVDA port map( A => n3337, Y => n4518, Z => n4706);
   U5132 : IVDA port map( A => n1475, Y => n_3426, Z => n4702);
   U5133 : IVDA port map( A => n1476, Y => n_3427, Z => n4701);
   U5134 : IVI port map( A => n4889, Z => n4888);
   U5135 : AO6 port map( A => n2650, B => n2651, C => n4379, Z => n2636);
   U5136 : NR4 port map( A => n2638, B => n2639, C => n2640, D => n2641, Z => 
                           n2637);
   U5137 : AO2 port map( A => v_RAM_OUT0_25_port, B => n2655, C => n5054, D => 
                           n5233, Z => n2650);
   U5138 : AO4 port map( A => n4552, B => n4404, C => v_RAM_OUT0_10_port, D => 
                           n2164, Z => n2160);
   U5139 : AO4 port map( A => n4766, B => n2162, C => n5134, D => n4413, Z => 
                           n2161);
   U5140 : AO4 port map( A => n4397, B => n2657, C => v_RAM_OUT0_26_port, D => 
                           n2658, Z => n2655);
   U5141 : AO2 port map( A => n2659, B => n1949, C => n5062, D => n4781, Z => 
                           n2658);
   U5142 : AO7 port map( A => v_RAM_OUT0_10_port, B => n2382, C => n2383, Z => 
                           n1892);
   U5143 : AO2 port map( A => n5144, B => n4769, C => n4766, D => n2320, Z => 
                           n2383);
   U5144 : AO2 port map( A => v_RAM_OUT0_12_port, B => n2384, C => n2298, D => 
                           n4404, Z => n2382);
   U5145 : AO3 port map( A => n1953, B => n4838, C => n2652, D => n2653, Z => 
                           n2651);
   U5146 : AO4 port map( A => n5055, B => n4727, C => n5064, D => n2505, Z => 
                           n2502);
   U5147 : AO6 port map( A => n5058, B => v_RAM_OUT0_26_port, C => n4839, Z => 
                           n2505);
   U5148 : AO3 port map( A => n3055, B => n2918, C => n3056, D => n4402, Z => 
                           n3045);
   U5149 : ND3 port map( A => n3057, B => n4395, C => v_RAM_OUT0_17_port, Z => 
                           n3056);
   U5150 : AO4 port map( A => n5079, B => n4715, C => n5089, D => n2912, Z => 
                           n2909);
   U5151 : AO6 port map( A => n5096, B => v_RAM_OUT0_18_port, C => n4356, Z => 
                           n2912);
   U5152 : AO4 port map( A => n5117, B => n4737, C => n2050, D => n2051, Z => 
                           n2047);
   U5153 : AO6 port map( A => n5133, B => v_RAM_OUT0_10_port, C => n4765, Z => 
                           n2051);
   U5154 : AO3 port map( A => n3458, B => n3321, C => n3459, D => n4401, Z => 
                           n3448);
   U5155 : ND3 port map( A => n3460, B => n4371, C => v_RAM_OUT0_1_port, Z => 
                           n3459);
   U5156 : AO4 port map( A => n5156, B => n4705, C => n5166, D => n3315, Z => 
                           n3312);
   U5157 : AO6 port map( A => n5173, B => v_RAM_OUT0_2_port, C => n4808, Z => 
                           n3315);
   U5158 : AO3 port map( A => n2070, B => n1884, C => n2387, D => n2388, Z => 
                           n2386);
   U5159 : EO1 port map( A => v_RAM_OUT0_25_port, B => n2877, C => n2612, D => 
                           n2511, Z => n2876);
   U5160 : AO3 port map( A => n4397, B => n2579, C => n5042, D => n2878, Z => 
                           n2877);
   U5161 : EO1 port map( A => n5041, B => n4781, C => n4828, D => n2647, Z => 
                           n2878);
   U5162 : AO2 port map( A => n4729, B => n2814, C => n2519, D => n1949, Z => 
                           n2813);
   U5163 : EO1 port map( A => v_RAM_OUT0_17_port, B => n3289, C => n3018, D => 
                           n2918, Z => n3288);
   U5164 : AO3 port map( A => n4395, B => n2986, C => n5085, D => n3290, Z => 
                           n3289);
   U5165 : EO1 port map( A => n5102, B => n4780, C => n4813, D => n3055, Z => 
                           n3290);
   U5166 : AO2 port map( A => n4716, B => n3202, C => n2927, D => n1696, Z => 
                           n3201);
   U5167 : EO1 port map( A => v_RAM_OUT0_1_port, B => n3697, C => n3421, D => 
                           n3321, Z => n3696);
   U5168 : AO3 port map( A => n4371, B => n3389, C => n5162, D => n3698, Z => 
                           n3697);
   U5169 : EO1 port map( A => n5179, B => n4779, C => n4797, D => n3458, Z => 
                           n3698);
   U5170 : AO2 port map( A => n4706, B => n3606, C => n3330, D => n2481, Z => 
                           n3605);
   U5171 : AO6 port map( A => n5131, B => v_RAM_OUT0_13_port, C => n2268, Z => 
                           n2315);
   U5172 : AO3 port map( A => n4416, B => n2511, C => n2835, D => n2836, Z => 
                           n2823);
   U5173 : AO2 port map( A => n5229, B => n2515, C => n5041, D => n5230, Z => 
                           n2836);
   U5174 : AO2 port map( A => n2837, B => n4729, C => n5063, D => n2519, Z => 
                           n2835);
   U5175 : AO7 port map( A => n2621, B => n2622, C => n5204, Z => n2620);
   U5176 : AO3 port map( A => n5029, B => n4828, C => n2623, D => n2618, Z => 
                           n2621);
   U5177 : AO4 port map( A => n1953, B => n4725, C => n4781, D => n2553, Z => 
                           n2622);
   U5178 : AO3 port map( A => n4399, B => n2918, C => n3240, D => n3241, Z => 
                           n3228);
   U5179 : AO2 port map( A => n5225, B => n2922, C => n5102, D => n5219, Z => 
                           n3241);
   U5180 : AO2 port map( A => n3242, B => n4716, C => n5088, D => n2927, Z => 
                           n3240);
   U5181 : AO7 port map( A => n3028, B => n3029, C => n5193, Z => n3027);
   U5182 : AO3 port map( A => n5107, B => n4813, C => n3030, D => n3024, Z => 
                           n3028);
   U5183 : AO4 port map( A => n1697, B => n4717, C => n4780, D => n2961, Z => 
                           n3029);
   U5184 : AO2 port map( A => n5070, B => n2088_port, C => n2089_port, D => 
                           n2090, Z => n2086_port);
   U5185 : AO6 port map( A => n5123, B => n4767, C => n4740, Z => n2089_port);
   U5186 : AO3 port map( A => n4739, B => n5125, C => n2097, D => n2098, Z => 
                           n2088_port);
   U5187 : AO4 port map( A => n5120, B => n2065, C => n2066, D => n2067, Z => 
                           n2063);
   U5188 : EON1 port map( A => n2070, B => n2071, C => n2046, D => n5203, Z => 
                           n2062);
   U5189 : AO3 port map( A => n4398, B => n3321, C => n3645, D => n3646, Z => 
                           n3633);
   U5190 : AO2 port map( A => n5216, B => n3325, C => n5179, D => n5210, Z => 
                           n3646);
   U5191 : AO2 port map( A => n3647, B => n4706, C => n5165, D => n3330, Z => 
                           n3645);
   U5192 : AO7 port map( A => n3431, B => n3432, C => n5206, Z => n3430);
   U5193 : AO3 port map( A => n5184, B => n4797, C => n3433, D => n3427, Z => 
                           n3431);
   U5194 : AO4 port map( A => n2482, B => n4707, C => n4779, D => n3364, Z => 
                           n3432);
   U5195 : AO7 port map( A => n4401, B => n2462, C => n2463, Z => n2461);
   U5196 : AO2 port map( A => n4522, B => n2464, C => n5163, D => n4386, Z => 
                           n2463);
   U5197 : AO4 port map( A => n5209, B => n2467, C => n2468, D => n2469, Z => 
                           n2464);
   U5198 : AO2 port map( A => v_RAM_OUT0_2_port, B => n2470, C => n5157, D => 
                           n4371, Z => n2468);
   U5199 : AO7 port map( A => v_RAM_OUT0_5_port, B => n2473, C => n2474, Z => 
                           n2460);
   U5200 : AO2 port map( A => n5207, B => n2476, C => n2477, D => n5206, Z => 
                           n2474);
   U5201 : AO4 port map( A => n5209, B => n2479, C => n2480, D => n2469, Z => 
                           n2476);
   U5202 : AO2 port map( A => v_RAM_OUT0_2_port, B => n2481, C => n2482, D => 
                           n4371, Z => n2480);
   U5203 : AO7 port map( A => n4379, B => n1958, C => n2864, Z => n2863);
   U5204 : AO2 port map( A => n4521, B => n2865, C => n5037, D => n4400, Z => 
                           n2864);
   U5205 : AO4 port map( A => n5227, B => n1962, C => n2871, D => n1954, Z => 
                           n2865);
   U5206 : AO2 port map( A => v_RAM_OUT0_26_port, B => n1964, C => n5049, D => 
                           n4397, Z => n2871);
   U5207 : AO7 port map( A => v_RAM_OUT0_29_port, B => n1946, C => n2879, Z => 
                           n2862);
   U5208 : AO2 port map( A => n5205, B => n2880, C => n1956, D => n5204, Z => 
                           n2879);
   U5209 : AO4 port map( A => n5227, B => n2532, C => n2883, D => n1954, Z => 
                           n2880);
   U5210 : AO2 port map( A => v_RAM_OUT0_26_port, B => n4724, C => n1953, D => 
                           n4397, Z => n2883);
   U5211 : AO7 port map( A => n4403, B => n1677, C => n1678, Z => n1676);
   U5212 : AO2 port map( A => n4520, B => n1679, C => n5086, D => n4385, Z => 
                           n1678);
   U5213 : AO4 port map( A => n5218, B => n1682, C => n1683, D => n1684, Z => 
                           n1679);
   U5214 : AO2 port map( A => v_RAM_OUT0_18_port, B => n1685, C => n5080, D => 
                           n4395, Z => n1683);
   U5215 : AO7 port map( A => n4782, B => n1688, C => n1689, Z => n1675);
   U5216 : AO2 port map( A => n5194, B => n1691, C => n1692, D => n5193, Z => 
                           n1689);
   U5217 : AO4 port map( A => n5218, B => n1694, C => n1695, D => n1684, Z => 
                           n1691);
   U5218 : AO2 port map( A => v_RAM_OUT0_18_port, B => n1696, C => n1697, D => 
                           n4395, Z => n1695);
   U5219 : AO4 port map( A => n1942, B => n4579, C => v_RAM_OUT0_31_port, D => 
                           n1943, Z => n1606);
   U5220 : AO2 port map( A => n1944, B => n1945, C => n1946, D => n4379, Z => 
                           n1943);
   U5221 : AO6 port map( A => v_RAM_OUT0_29_port, B => n1958, C => n1959, Z => 
                           n1942);
   U5222 : AO6 port map( A => n1956, B => n4510, C => n4379, Z => n1944);
   U5223 : AO7 port map( A => v_RAM_OUT0_31_port, B => n2821, C => n2822, Z => 
                           n1601);
   U5224 : AO6 port map( A => v_RAM_OUT0_29_port, B => n2838, C => n2839, Z => 
                           n2821);
   U5225 : AO3 port map( A => n2823, B => n2824, C => v_RAM_OUT0_31_port, D => 
                           n2825, Z => n2822);
   U5226 : ND4 port map( A => n2850, B => n2851, C => n2852, D => n2853, Z => 
                           n2838);
   U5227 : AO4 port map( A => v_RAM_OUT0_31_port, B => n5030, C => n1917, D => 
                           n4579, Z => n1595);
   U5228 : AO6 port map( A => v_RAM_OUT0_29_port, B => n1919, C => n1920, Z => 
                           n1917);
   U5229 : AO4 port map( A => n5028, B => n4730, C => n1923, D => n4731, Z => 
                           n1920);
   U5230 : AO7 port map( A => v_RAM_OUT0_31_port, B => n2739, C => n2740, Z => 
                           n1590);
   U5231 : AO6 port map( A => v_RAM_OUT0_29_port, B => n2762, C => n2763, Z => 
                           n2739);
   U5232 : AO3 port map( A => n2741, B => n2742, C => v_RAM_OUT0_31_port, D => 
                           n2743, Z => n2740);
   U5233 : AO4 port map( A => n2764, B => n4731, C => n2765, D => n4730, Z => 
                           n2763);
   U5234 : AO4 port map( A => n3265, B => n4564, C => v_RAM_OUT0_23_port, D => 
                           n3266, Z => n1813);
   U5235 : AO2 port map( A => n3267, B => n3268, C => n1688, D => n4402, Z => 
                           n3266);
   U5236 : AO6 port map( A => n4782, B => n1677, C => n3277, Z => n3265);
   U5237 : AO6 port map( A => n1692, B => n4509, C => n4403, Z => n3267);
   U5238 : AO7 port map( A => v_RAM_OUT0_23_port, B => n3226, C => n3227, Z => 
                           n1663);
   U5239 : AO6 port map( A => n4782, B => n3243, C => n3244, Z => n3226);
   U5240 : AO3 port map( A => n3228, B => n3229, C => v_RAM_OUT0_23_port, D => 
                           n3230, Z => n3227);
   U5241 : ND4 port map( A => n3255, B => n3256, C => n3257, D => n3258, Z => 
                           n3243);
   U5242 : AO4 port map( A => v_RAM_OUT0_23_port, B => n5084, C => n3190, D => 
                           n4564, Z => n1805);
   U5243 : AO6 port map( A => n4782, B => n1648, C => n3191, Z => n3190);
   U5244 : AO4 port map( A => n5092, B => n4721, C => n3192, D => n4720, Z => 
                           n3191);
   U5245 : AO7 port map( A => v_RAM_OUT0_23_port, B => n3146, C => n3147, Z => 
                           n1632);
   U5246 : AO6 port map( A => n4782, B => n3169, C => n3170, Z => n3146);
   U5247 : AO3 port map( A => n3148, B => n3149, C => v_RAM_OUT0_23_port, D => 
                           n3150, Z => n3147);
   U5248 : AO4 port map( A => n3171, B => n4720, C => n3172, D => n4721, Z => 
                           n3170);
   U5249 : AO4 port map( A => n3673, B => n4580, C => v_RAM_OUT0_7_port, D => 
                           n3674, Z => n1562);
   U5250 : AO2 port map( A => n3675, B => n3676, C => n2473, D => n4401, Z => 
                           n3674);
   U5251 : AO6 port map( A => v_RAM_OUT0_5_port, B => n2462, C => n3685, Z => 
                           n3673);
   U5252 : AO6 port map( A => n2477, B => n4508, C => n4401, Z => n3675);
   U5253 : AO7 port map( A => v_RAM_OUT0_7_port, B => n3631, C => n3632, Z => 
                           n1557);
   U5254 : AO6 port map( A => v_RAM_OUT0_5_port, B => n3648, C => n3649, Z => 
                           n3631);
   U5255 : AO3 port map( A => n3633, B => n3634, C => v_RAM_OUT0_7_port, D => 
                           n3635, Z => n3632);
   U5256 : ND4 port map( A => n3660, B => n3661, C => n3662, D => n3663, Z => 
                           n3648);
   U5257 : AO4 port map( A => v_RAM_OUT0_7_port, B => n5161, C => n3594, D => 
                           n4580, Z => n1551);
   U5258 : AO6 port map( A => v_RAM_OUT0_5_port, B => n2437, C => n3595, Z => 
                           n3594);
   U5259 : AO4 port map( A => n5169, B => n4711, C => n3596, D => n4710, Z => 
                           n3595);
   U5260 : AO7 port map( A => v_RAM_OUT0_7_port, B => n3550, C => n3551, Z => 
                           n1545);
   U5261 : AO6 port map( A => v_RAM_OUT0_5_port, B => n3573, C => n3574, Z => 
                           n3550);
   U5262 : AO3 port map( A => n3552, B => n3553, C => v_RAM_OUT0_7_port, D => 
                           n3554, Z => n3551);
   U5263 : AO4 port map( A => n3575, B => n4710, C => n3576, D => n4711, Z => 
                           n3574);
   U5264 : AO6 port map( A => n5226, B => n2575, C => n5228, Z => n2776);
   U5265 : AO6 port map( A => n5217, B => n2982, C => n5224, Z => n3183);
   U5266 : AO6 port map( A => n5208, B => n3385, C => n5215, Z => n3587);
   U5267 : AO4 port map( A => n2633, B => n2634, C => v_RAM_OUT0_31_port, D => 
                           n2635, Z => n2632);
   U5268 : AO3 port map( A => n2671, B => n4730, C => n2672, D => n5040, Z => 
                           n2633);
   U5269 : AO3 port map( A => n1606, B => n1758, C => n1784, D => n1785, Z => 
                           n4257);
   U5270 : AO7 port map( A => n4685, B => n4855, C => n4752, Z => n1786);
   U5271 : AO3 port map( A => n1590, B => n1758, C => n1773, D => n1774, Z => 
                           n4260);
   U5272 : AO7 port map( A => n4688, B => n4855, C => n4751, Z => n1775);
   U5273 : AO3 port map( A => n5033, B => n1758, C => n1766, D => n1767, Z => 
                           n4262);
   U5274 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n4855, C => n4751, Z 
                           => n1768);
   U5275 : AO3 port map( A => n1663, B => n1787, C => n1810, D => n1811, Z => 
                           n4266);
   U5276 : AO7 port map( A => n4679, B => n4856, C => n4749, Z => n1812);
   U5277 : AO3 port map( A => n1628, B => n1787, C => n1798, D => n1799, Z => 
                           n4269);
   U5278 : AO7 port map( A => v_KEY_COLUMN_20_port, B => n4855, C => n4750, Z 
                           => n1800);
   U5279 : AO3 port map( A => n5065, B => n1787, C => n1795, D => n1796, Z => 
                           n4270);
   U5280 : AO7 port map( A => n4682, B => n4855, C => n4749, Z => n1797);
   U5281 : AO3 port map( A => n1836, B => n1818, C => n1837, D => n1838, Z => 
                           n4275);
   U5282 : AO6 port map( A => n5066, B => v_RAM_OUT0_9_port, C => n1841, Z => 
                           n1836);
   U5283 : AO3 port map( A => n1498, B => n1818, C => n1830, D => n1831, Z => 
                           n4277);
   U5284 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n4856, C => n4748, Z 
                           => n1832);
   U5285 : AO3 port map( A => n1562, B => n3291, C => n3667, D => n3668, Z => 
                           n4281);
   U5286 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n4855, C => n4713, Z =>
                           n3670);
   U5287 : AO3 port map( A => n1557, B => n3291, C => n3627, D => n3628, Z => 
                           n4282);
   U5288 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n4856, C => n4712, Z =>
                           n3630);
   U5289 : AO3 port map( A => n1551, B => n3291, C => n3590, D => n3591, Z => 
                           n4283);
   U5290 : AO7 port map( A => n4669, B => n4855, C => n4713, Z => n3593);
   U5291 : AO3 port map( A => n1545, B => n3291, C => n3546, D => n3547, Z => 
                           n4284);
   U5292 : AO7 port map( A => n4670, B => n4856, C => n4712, Z => n3549);
   U5293 : AO3 port map( A => n1539, B => n3291, C => n3500, D => n3501, Z => 
                           n4285);
   U5294 : AO7 port map( A => n4671, B => n4856, C => n4713, Z => n3503);
   U5295 : AO3 port map( A => n5073, B => n3291, C => n3439, D => n3440, Z => 
                           n4286);
   U5296 : AO7 port map( A => v_KEY_COLUMN_5_port, B => n4856, C => n4712, Z =>
                           n3441);
   U5297 : EON1 port map( A => n4369, B => n1413, C => N2085, D => n1409, Z => 
                           n4310);
   U5298 : ND4 port map( A => n2992, B => n2993, C => n2994, D => n2995, Z => 
                           n2973);
   U5299 : AO2 port map( A => n5112, B => n5221, C => n5225, D => n3003, Z => 
                           n2994);
   U5300 : AO2 port map( A => n5222, B => n3007, C => n2964, D => n5224, Z => 
                           n2992);
   U5301 : AO2 port map( A => n2996, B => v_RAM_OUT0_17_port, C => n5107, D => 
                           n4509, Z => n2995);
   U5302 : NR4 port map( A => n2248, B => n2249, C => n5199, D => n2250, Z => 
                           n2233);
   U5303 : NR3 port map( A => n2033, B => v_RAM_OUT0_13_port, C => 
                           v_RAM_OUT0_12_port, Z => n2249);
   U5304 : AO4 port map( A => n4736, B => n2073, C => n2251, D => n1857, Z => 
                           n2248);
   U5305 : AO3 port map( A => n2391, B => n4739, C => n2392, D => n2393, Z => 
                           n1873);
   U5306 : AO7 port map( A => n2394, B => n5145, C => v_RAM_OUT0_10_port, Z => 
                           n2392);
   U5307 : AO2 port map( A => n4504, B => n2094, C => n4767, D => n2200, Z => 
                           n2393);
   U5308 : ND4 port map( A => n2715, B => n2716, C => n2717, D => n2718, Z => 
                           n2693);
   U5309 : ND4 port map( A => n2695, B => v_RAM_OUT0_31_port, C => n2696, D => 
                           n2697, Z => n2694);
   U5310 : AO7 port map( A => n2719, B => n2720, C => n5205, Z => n2718);
   U5311 : ND4 port map( A => n3121, B => n3122, C => n3123, D => n3124, Z => 
                           n3100);
   U5312 : ND4 port map( A => n3102, B => v_RAM_OUT0_23_port, C => n3103, D => 
                           n3104, Z => n3101);
   U5313 : AO7 port map( A => n3125, B => n3126, C => n5194, Z => n3124);
   U5314 : ND4 port map( A => n3525, B => n3526, C => n3527, D => n3528, Z => 
                           n3504);
   U5315 : ND4 port map( A => n3506, B => v_RAM_OUT0_7_port, C => n3507, D => 
                           n3508, Z => n3505);
   U5316 : AO7 port map( A => n3529, B => n3530, C => n5207, Z => n3528);
   U5317 : IVDA port map( A => n1472, Y => n4428, Z => n4697);
   U5318 : AO4 port map( A => n4731, B => n2544, C => n4730, D => n4724, Z => 
                           n2539);
   U5319 : AO4 port map( A => n4720, B => n2951, C => n4721, D => n1696, Z => 
                           n2947);
   U5320 : AO4 port map( A => n4710, B => n3354, C => n4711, D => n2481, Z => 
                           n3350);
   U5321 : ND4 port map( A => n2884, B => n2885, C => n2886, D => n2887, Z => 
                           n1946);
   U5322 : AO2 port map( A => n5229, B => n4416, C => n5228, D => n2815, Z => 
                           n2884);
   U5323 : AO2 port map( A => n5076, B => n5232, C => n4729, D => n2610, Z => 
                           n2887);
   U5324 : ND4 port map( A => n3269, B => n3270, C => n3271, D => n3272, Z => 
                           n1688);
   U5325 : AO2 port map( A => n5225, B => n4399, C => n5224, D => n3204, Z => 
                           n3269);
   U5326 : AO2 port map( A => n5087, B => n5221, C => n4716, D => n3016, Z => 
                           n3272);
   U5327 : ND4 port map( A => n3677, B => n3678, C => n3679, D => n3680, Z => 
                           n2473);
   U5328 : AO2 port map( A => n5216, B => n4398, C => n5215, D => n3608, Z => 
                           n3677);
   U5329 : AO2 port map( A => n5164, B => n5212, C => n4706, D => n3419, Z => 
                           n3680);
   U5330 : AO6 port map( A => n2961, B => n3077, C => n4823, Z => n3074);
   U5331 : AO6 port map( A => n3364, B => n3480, C => n4807, Z => n3477);
   U5332 : AO3 port map( A => n2647, B => n2511, C => n2648, D => n4379, Z => 
                           n2638);
   U5333 : ND3 port map( A => n2649, B => n4397, C => v_RAM_OUT0_25_port, Z => 
                           n2648);
   U5334 : AO6 port map( A => n2094, B => n2095, C => n4412, Z => n2091);
   U5335 : NR3 port map( A => n5046, B => n2881, C => n2882, Z => n1956);
   U5336 : AO4 port map( A => n4827, B => n4724, C => n5057, D => n4837, Z => 
                           n2881);
   U5337 : AO4 port map( A => n4781, B => n2520, C => n2645, D => n1966, Z => 
                           n2882);
   U5338 : NR3 port map( A => n5236, B => n3275, C => n3276, Z => n1692);
   U5339 : AO4 port map( A => n4812, B => n4719, C => n5112, D => n4822, Z => 
                           n3275);
   U5340 : AO4 port map( A => n4780, B => n2928, C => n3052, D => n4714, Z => 
                           n3276);
   U5341 : AO2 port map( A => n2010, B => v_RAM_OUT0_13_port, C => n5195, D => 
                           n2012, Z => n2009);
   U5342 : NR3 port map( A => n5243, B => n3683, C => n3684, Z => n2477);
   U5343 : AO4 port map( A => n4796, B => n4709, C => n5189, D => n4806, Z => 
                           n3683);
   U5344 : AO4 port map( A => n4779, B => n3331, C => n3455, D => n4704, Z => 
                           n3684);
   U5345 : AO3 port map( A => n5076, B => n2578, C => v_RAM_OUT0_29_port, D => 
                           n2833, Z => n2824);
   U5346 : EO1 port map( A => n2647, B => n5226, C => n2522, D => n1931, Z => 
                           n2833);
   U5347 : AO2 port map( A => n5204, B => n2710, C => n4400, D => n2711, Z => 
                           n2695);
   U5348 : AO3 port map( A => v_RAM_OUT0_26_port, B => n2553, C => n5038, D => 
                           n2713, Z => n2710);
   U5349 : AO3 port map( A => n4726, B => n2700, C => n4827, D => n2712, Z => 
                           n2711);
   U5350 : AO2 port map( A => n5045, B => n5231, C => n4839, D => n2714, Z => 
                           n2713);
   U5351 : AO3 port map( A => n5087, B => n2985, C => n4782, D => n3238, Z => 
                           n3229);
   U5352 : EO1 port map( A => n3055, B => n5217, C => n2931, D => n1658, Z => 
                           n3238);
   U5353 : AO3 port map( A => n3159, B => n3051, C => n4782, D => n3160, Z => 
                           n3149);
   U5354 : AO2 port map( A => n5221, B => n2966, C => n5217, D => n3161, Z => 
                           n3160);
   U5355 : AO2 port map( A => n5193, B => n3116, C => n4385, D => n3117, Z => 
                           n3102);
   U5356 : AO3 port map( A => v_RAM_OUT0_18_port, B => n2961, C => n5093, D => 
                           n3119, Z => n3116);
   U5357 : AO3 port map( A => n4718, B => n3107, C => n4812, D => n3118, Z => 
                           n3117);
   U5358 : AO2 port map( A => n5115, B => n5220, C => n4356, D => n3120, Z => 
                           n3119);
   U5359 : AO3 port map( A => n5164, B => n3388, C => v_RAM_OUT0_5_port, D => 
                           n3643, Z => n3634);
   U5360 : EO1 port map( A => n3458, B => n5208, C => n3334, D => n2447, Z => 
                           n3643);
   U5361 : AO3 port map( A => n3563, B => n3454, C => v_RAM_OUT0_5_port, D => 
                           n3564, Z => n3553);
   U5362 : AO2 port map( A => n5212, B => n3369, C => n5208, D => n3565, Z => 
                           n3564);
   U5363 : AO2 port map( A => n5206, B => n3520, C => n4386, D => n3521, Z => 
                           n3506);
   U5364 : AO3 port map( A => v_RAM_OUT0_2_port, B => n3364, C => n5170, D => 
                           n3523, Z => n3520);
   U5365 : AO3 port map( A => n4708, B => n3511, C => n4796, D => n3522, Z => 
                           n3521);
   U5366 : AO2 port map( A => n5192, B => n5211, C => n4808, D => n3524, Z => 
                           n3523);
   U5367 : AO7 port map( A => n4401, B => n2437, C => n2438, Z => n2433);
   U5368 : AO2 port map( A => n5169, B => n4522, C => n4386, D => n2442, Z => 
                           n2438);
   U5369 : AO2 port map( A => n5181, B => n5214, C => n5191, D => 
                           v_RAM_OUT0_2_port, Z => n2443);
   U5370 : AO7 port map( A => n4379, B => n1919, C => n2802, Z => n2784);
   U5371 : AO2 port map( A => n5028, B => n4521, C => n4400, D => n2803, Z => 
                           n2802);
   U5372 : AO2 port map( A => n5044, B => n5234, C => n5060, D => 
                           v_RAM_OUT0_26_port, Z => n2804);
   U5373 : AO7 port map( A => n4402, B => n1648, C => n1649, Z => n1644);
   U5374 : AO2 port map( A => n5092, B => n4520, C => n4385, D => n1653, Z => 
                           n1649);
   U5375 : AO2 port map( A => n5104, B => n5223, C => n5114, D => 
                           v_RAM_OUT0_18_port, Z => n1654);
   U5376 : AO3 port map( A => n1954, B => n2668, C => n2807, D => n2808, Z => 
                           n2806);
   U5377 : AO2 port map( A => n5036, B => n5231, C => n5029, D => n5234, Z => 
                           n2808);
   U5378 : AO3 port map( A => n1684, B => n3076, C => n3196, D => n3197, Z => 
                           n3195);
   U5379 : AO2 port map( A => n5111, B => n5220, C => n5107, D => n5223, Z => 
                           n3197);
   U5380 : AO3 port map( A => n2469, B => n3479, C => n3600, D => n3601, Z => 
                           n3599);
   U5381 : AO2 port map( A => n5188, B => n5211, C => n5184, D => n5214, Z => 
                           n3601);
   U5382 : AO3 port map( A => n4823, B => n3018, C => n4385, D => n3019, Z => 
                           n3008);
   U5383 : AO6 port map( A => n3023, B => n3024, C => n4715, Z => n3022);
   U5384 : AO3 port map( A => n5087, B => n4823, C => n4520, D => n3010, Z => 
                           n3009);
   U5385 : AO6 port map( A => n3015, B => n3016, C => n4718, Z => n3013);
   U5386 : AO3 port map( A => n2210, B => n2173, C => n2211, D => n2212, Z => 
                           n2209);
   U5387 : AO7 port map( A => n2213, B => n5198, C => n2214, Z => n2212);
   U5388 : ND4 port map( A => n2586, B => n2587, C => n2588, D => n2589, Z => 
                           n2567);
   U5389 : AO2 port map( A => n5057, B => n5232, C => n5229, D => n1930, Z => 
                           n2588);
   U5390 : AO2 port map( A => n5233, B => n2600, C => n2556, D => n5228, Z => 
                           n2586);
   U5391 : AO2 port map( A => n2590, B => v_RAM_OUT0_25_port, C => n5029, D => 
                           n4510, Z => n2589);
   U5392 : ND4 port map( A => n3395, B => n3396, C => n3397, D => n3398, Z => 
                           n3376);
   U5393 : AO2 port map( A => n5189, B => n5212, C => n5216, D => n3406, Z => 
                           n3397);
   U5394 : AO2 port map( A => n5213, B => n3410, C => n3367, D => n5215, Z => 
                           n3395);
   U5395 : AO2 port map( A => n3399, B => v_RAM_OUT0_1_port, C => n5184, D => 
                           n4508, Z => n3398);
   U5396 : AO2 port map( A => n5123, B => n4515, C => n4768, D => n2298, Z => 
                           n2401);
   U5397 : AO2 port map( A => n4504, B => n2094, C => n4765, D => n4405, Z => 
                           n2402);
   U5398 : AO6 port map( A => n2162, B => n2164, C => n4738, Z => n2338);
   U5399 : AO7 port map( A => v_RAM_OUT0_24_port, B => n4837, C => n4727, Z => 
                           n1926);
   U5400 : AO7 port map( A => v_RAM_OUT0_16_port, B => n4822, C => n4714, Z => 
                           n1656);
   U5401 : AO7 port map( A => v_RAM_OUT0_0_port, B => n4806, C => n4704, Z => 
                           n2445);
   U5402 : IVDA port map( A => n1922, Y => n4521, Z => n4730);
   U5403 : IVDA port map( A => n2901, Y => n4520, Z => n4721);
   U5404 : IVDA port map( A => n3304, Y => n4522, Z => n4711);
   U5405 : IVDA port map( A => n1469, Y => n_3428, Z => n4699);
   U5406 : IVDA port map( A => n1470, Y => n_3429, Z => n4698);
   U5407 : IVDA port map( A => n1465, Y => n_3430, Z => n4695);
   U5408 : AO6 port map( A => n2731, B => n2732, C => n4827, Z => n2729);
   U5409 : AO6 port map( A => n3137, B => n3138, C => n4812, Z => n3135);
   U5410 : AO6 port map( A => n3541, B => n3542, C => n4796, Z => n3539);
   U5411 : AO2 port map( A => n4695, B => n4590, C => n4696, D => n4432, Z => 
                           n3793);
   U5412 : AO2 port map( A => n4693, B => n4433, C => n4694, D => n4595, Z => 
                           n3792);
   U5413 : AO2 port map( A => n4695, B => n4591, C => n4696, D => n4467, Z => 
                           n3782);
   U5414 : AO2 port map( A => n4693, B => n4434, C => n4694, D => n4596, Z => 
                           n3781);
   U5415 : AO2 port map( A => n4695, B => n4592, C => n4696, D => n4468, Z => 
                           n3771);
   U5416 : AO2 port map( A => n4693, B => n4435, C => n4694, D => n4383, Z => 
                           n3770);
   U5417 : AO2 port map( A => n4695, B => n4593, C => n4696, D => n4441, Z => 
                           n3760);
   U5418 : AO2 port map( A => n4693, B => n4388, C => n4694, D => n4444, Z => 
                           n3759);
   U5419 : AO2 port map( A => n4695, B => n4594, C => n4696, D => n4469, Z => 
                           n3749);
   U5420 : AO2 port map( A => n4693, B => n4557, C => n4694, D => n4445, Z => 
                           n3748);
   U5421 : AO2 port map( A => n4695, B => n4409, C => n4696, D => n4529, Z => 
                           n3738);
   U5422 : AO2 port map( A => n4693, B => n4470, C => n4694, D => n4597, Z => 
                           n3737);
   U5423 : AO2 port map( A => n4695, B => n4524, C => n4696, D => n4417, Z => 
                           n3726);
   U5424 : AO2 port map( A => n4693, B => n4382, C => n4694, D => n4421, Z => 
                           n3725);
   U5425 : AO2 port map( A => n4695, B => n4438, C => n4696, D => n4530, Z => 
                           n3713);
   U5426 : AO2 port map( A => n4693, B => n4531, C => n4694, D => n4410, Z => 
                           n3712);
   U5427 : AO3 port map( A => n2752, B => n2644, C => v_RAM_OUT0_29_port, D => 
                           n2753, Z => n2742);
   U5428 : AO2 port map( A => n5232, B => n2559, C => n5226, D => n2754, Z => 
                           n2753);
   U5429 : AO2 port map( A => n2703, B => n2683, C => n4521, D => n2704, Z => 
                           n2696);
   U5430 : AO4 port map( A => n4838, B => n2677, C => n5060, D => n2706, Z => 
                           n2704);
   U5431 : AO6 port map( A => n5034, B => n4781, C => n5231, Z => n2706);
   U5432 : AO6 port map( A => n5204, B => n2723, C => v_RAM_OUT0_31_port, Z => 
                           n2717);
   U5433 : AO3 port map( A => n4725, B => n2541, C => n2724, D => n2725, Z => 
                           n2723);
   U5434 : AO7 port map( A => n5051, B => n5059, C => n4831, Z => n2724);
   U5435 : AO2 port map( A => n5064, B => n5231, C => n4839, D => n2612, Z => 
                           n2725);
   U5436 : AO3 port map( A => n4837, B => n2646, C => n4521, D => n2727, Z => 
                           n2716);
   U5437 : AO6 port map( A => n2575, B => n2574, C => n4726, Z => n2730);
   U5438 : AO2 port map( A => n3110, B => n3091, C => n4520, D => n3111, Z => 
                           n3103);
   U5439 : AO4 port map( A => n4823, B => n3085, C => n5114, D => n3112, Z => 
                           n3111);
   U5440 : AO6 port map( A => n5109, B => n4780, C => n5220, Z => n3112);
   U5441 : AO6 port map( A => n5193, B => n3129, C => v_RAM_OUT0_23_port, Z => 
                           n3123);
   U5442 : AO3 port map( A => n4717, B => n2949, C => n3130, D => n3131, Z => 
                           n3129);
   U5443 : AO7 port map( A => n5090, B => n5237, C => n4816, Z => n3130);
   U5444 : AO2 port map( A => n5089, B => n5220, C => n4356, D => n3018, Z => 
                           n3131);
   U5445 : AO3 port map( A => n4823, B => n3053, C => n4520, D => n3133, Z => 
                           n3122);
   U5446 : AO6 port map( A => n2982, B => n2981, C => n4718, Z => n3136);
   U5447 : AO3 port map( A => n4377, B => n1884, C => n2243, D => n2244, Z => 
                           n2234);
   U5448 : AO6 port map( A => n5148, B => n4767, C => n4740, Z => n2244);
   U5449 : AO2 port map( A => n4515, B => n2246, C => n2055, D => n4504, Z => 
                           n2243);
   U5450 : AO7 port map( A => n4776, B => n4405, C => n2068, Z => n2246);
   U5451 : AO2 port map( A => n3514, B => n3494, C => n4522, D => n3515, Z => 
                           n3507);
   U5452 : AO4 port map( A => n4807, B => n3488, C => n5191, D => n3516, Z => 
                           n3515);
   U5453 : AO6 port map( A => n5186, B => n4779, C => n5211, Z => n3516);
   U5454 : AO6 port map( A => n5206, B => n3533, C => v_RAM_OUT0_7_port, Z => 
                           n3527);
   U5455 : AO3 port map( A => n4707, B => n3352, C => n3534, D => n3535, Z => 
                           n3533);
   U5456 : AO7 port map( A => n5167, B => n5244, C => n4800, Z => n3534);
   U5457 : AO2 port map( A => n5166, B => n5211, C => n4808, D => n3421, Z => 
                           n3535);
   U5458 : AO3 port map( A => n4807, B => n3456, C => n4522, D => n3537, Z => 
                           n3526);
   U5459 : AO6 port map( A => n3385, B => n3384, C => n4708, Z => n3540);
   U5460 : AO3 port map( A => n5076, B => n4838, C => n4521, D => n2604, Z => 
                           n2602);
   U5461 : AO6 port map( A => n2609, B => n2610, C => n4726, Z => n2607);
   U5462 : AO3 port map( A => n4838, B => n2612, C => n4400, D => n2613, Z => 
                           n2601);
   U5463 : AO6 port map( A => n2617, B => n2618, C => n4727, Z => n2616);
   U5464 : AO3 port map( A => n5164, B => n4807, C => n4522, D => n3413, Z => 
                           n3412);
   U5465 : AO6 port map( A => n3418, B => n3419, C => n4708, Z => n3416);
   U5466 : AO3 port map( A => n4807, B => n3421, C => n4386, D => n3422, Z => 
                           n3411);
   U5467 : AO6 port map( A => n3426, B => n3427, C => n4705, Z => n3425);
   U5468 : AO6 port map( A => n2553, B => n2669, C => n4838, Z => n2666);
   U5469 : AO4 port map( A => n4728, B => n2609, C => n2722, D => n4837, Z => 
                           n2719);
   U5470 : AO4 port map( A => n4714, B => n3015, C => n3128, D => n4823, Z => 
                           n3125);
   U5471 : AO4 port map( A => n4704, B => n3418, C => n3532, D => n4807, Z => 
                           n3529);
   U5472 : AO4 port map( A => n4472, B => n4867, C => n4868, D => n4634, Z => 
                           n3970);
   U5473 : AO4 port map( A => n4473, B => n4866, C => n4871, D => n4635, Z => 
                           n3976);
   U5474 : AO4 port map( A => n4474, B => n4865, C => n4883, D => n4636, Z => 
                           n3982);
   U5475 : AO4 port map( A => n4475, B => n4865, C => n4880, D => n4637, Z => 
                           n3988);
   U5476 : AO4 port map( A => n4476, B => n4867, C => n4869, D => n4638, Z => 
                           n3994);
   U5477 : AO4 port map( A => n4477, B => n4866, C => n4873, D => n4639, Z => 
                           n4000);
   U5478 : AO4 port map( A => n4478, B => n4865, C => n4877, D => n4640, Z => 
                           n4006);
   U5479 : AO4 port map( A => n4479, B => n4867, C => n4868, D => n4641, Z => 
                           n4012);
   U5480 : AO4 port map( A => n4480, B => n4865, C => n4877, D => n4642, Z => 
                           n4018);
   U5481 : AO4 port map( A => n4481, B => n4866, C => n4872, D => n4643, Z => 
                           n4024);
   U5482 : AO4 port map( A => n4482, B => n4866, C => n4876, D => n4644, Z => 
                           n4030);
   U5483 : AO4 port map( A => n4483, B => n4866, C => n4873, D => n4645, Z => 
                           n4037);
   U5484 : AO4 port map( A => n4484, B => n4865, C => n4881, D => n4646, Z => 
                           n4043);
   U5485 : AO4 port map( A => n4485, B => n4866, C => n4874, D => n4647, Z => 
                           n4049);
   U5486 : AO4 port map( A => n4486, B => n4867, C => n4869, D => n4648, Z => 
                           n4055);
   U5487 : AO4 port map( A => n4487, B => n4865, C => n4878, D => n4649, Z => 
                           n4061);
   U5488 : AO4 port map( A => n4488, B => n4865, C => n4883, D => n4650, Z => 
                           n4067);
   U5489 : AO4 port map( A => n4489, B => n4866, C => n4872, D => n4651, Z => 
                           n4073);
   U5490 : AO4 port map( A => n4490, B => n4865, C => n4879, D => n4652, Z => 
                           n4080);
   U5491 : AO4 port map( A => n4491, B => n4865, C => n4881, D => n4653, Z => 
                           n4086);
   U5492 : AO4 port map( A => n4492, B => n4865, C => n4878, D => n4654, Z => 
                           n4092);
   U5493 : AO4 port map( A => n4493, B => n4866, C => n4870, D => n4655, Z => 
                           n4098);
   U5494 : AO4 port map( A => n4494, B => n4866, C => n4874, D => n4656, Z => 
                           n4104);
   U5495 : AO4 port map( A => n4495, B => n4865, C => n4882, D => n4657, Z => 
                           n4111);
   U5496 : AO4 port map( A => n4496, B => n4866, C => n4870, D => n4658, Z => 
                           n4117);
   U5497 : AO4 port map( A => n4497, B => n4866, C => n4875, D => n4659, Z => 
                           n4123);
   U5498 : AO4 port map( A => n4498, B => n4865, C => n4879, D => n4660, Z => 
                           n4129);
   U5499 : AO4 port map( A => n4499, B => n4865, C => n4882, D => n4661, Z => 
                           n4136);
   U5500 : AO4 port map( A => n4500, B => n4866, C => n4871, D => n4662, Z => 
                           n4142);
   U5501 : AO4 port map( A => n4501, B => n4866, C => n4875, D => n4663, Z => 
                           n4148);
   U5502 : AO4 port map( A => n4502, B => n4865, C => n4880, D => n4664, Z => 
                           n4154);
   U5503 : AO4 port map( A => n4503, B => n4866, C => n4876, D => n4665, Z => 
                           n4161);
   U5504 : AO3 port map( A => n4466, B => n1426, C => n5002, D => n4867, Z => 
                           n1445);
   U5505 : AO7 port map( A => n5027, B => n4604, C => n1457, Z => n1450);
   U5506 : AO7 port map( A => n4892, B => n1360, C => n5010, Z => n1446);
   U5507 : ND3 port map( A => n5010, B => n4603, C => n1452, Z => n1453);
   U5508 : ND4 port map( A => n5014, B => n1450, C => n4556, D => n4369, Z => 
                           n1454);
   U5509 : ND3 port map( A => n5010, B => n4366, C => n1452, Z => n1448);
   U5510 : AO3 port map( A => n4890, B => n4363, C => n1450, D => n1451, Z => 
                           n1449);
   U5511 : IVDA port map( A => n1388, Y => n4464, Z => n4703);
   U5512 : IVDA port map( A => n1370, Y => n4463, Z => n4762);
   U5513 : AO4 port map( A => n4463, B => n4600, C => n4998, D => n4762, Z => 
                           n4323);
   U5514 : AO4 port map( A => n4464, B => n4601, C => n4998, D => n4703, Z => 
                           n4331);
   U5515 : AO4 port map( A => n4465, B => n4602, C => n4761, D => n4998, Z => 
                           n4339);
   U5516 : AO7 port map( A => n1348, B => n4892, C => n5010, Z => n105);
   U5517 : AO6 port map( A => n3958, B => n1349, C => n1301, Z => n1348);
   U5518 : NR3 port map( A => v_CALCULATION_CNTR_0_port, B => 
                           v_CALCULATION_CNTR_3_port, C => n1457, Z => n3671);
   U5519 : AO3 port map( A => n4887, B => n4478, C => n522, D => n523, Z => 
                           n4010);
   U5520 : AO2 port map( A => n4784, B => n550, C => n551, D => n4787, Z => 
                           n522);
   U5521 : AO6 port map( A => n524, B => n4790, C => n525, Z => n523);
   U5522 : AO3 port map( A => n4888, B => n4491, C => n266, D => n267, Z => 
                           n4090);
   U5523 : AO2 port map( A => n4784, B => n290, C => n291, D => n4787, Z => 
                           n266);
   U5524 : AO6 port map( A => n268, B => n4790, C => n269, Z => n267);
   U5525 : AO3 port map( A => n4887, B => n4492, C => n464, D => n465, Z => 
                           n4096);
   U5526 : AO2 port map( A => n4784, B => n488, C => n489, D => n4787, Z => 
                           n464);
   U5527 : AO6 port map( A => n466, B => n4790, C => n467, Z => n465);
   U5528 : AO3 port map( A => n4888, B => n4475, C => n332, D => n333, Z => 
                           n3992);
   U5529 : AO2 port map( A => n4784, B => n362, C => n363, D => n4787, Z => 
                           n332);
   U5530 : AO6 port map( A => n334, B => n4790, C => n335, Z => n333);
   U5531 : AO3 port map( A => n4886, B => n4476, C => n1160, D => n1161, Z => 
                           n3998);
   U5532 : AO2 port map( A => n4783, B => n1200, C => n1201, D => n4788, Z => 
                           n1160);
   U5533 : AO6 port map( A => n1162, B => n4789, C => n1163, Z => n1161);
   U5534 : AO3 port map( A => n4887, B => n4477, C => n834, D => n835, Z => 
                           n4004);
   U5535 : AO2 port map( A => n4783, B => n873, C => n874, D => n4788, Z => 
                           n834);
   U5536 : AO6 port map( A => n836, B => n4789, C => n837, Z => n835);
   U5537 : AO3 port map( A => n4887, B => n4480, C => n561, D => n562, Z => 
                           n4022);
   U5538 : AO2 port map( A => n4784, B => n585, C => n586, D => n4787, Z => 
                           n561);
   U5539 : AO6 port map( A => n563, B => n4790, C => n564, Z => n562);
   U5540 : AO3 port map( A => n4886, B => n4481, C => n928, D => n929, Z => 
                           n4028);
   U5541 : AO2 port map( A => n4783, B => n959, C => n960, D => n4788, Z => 
                           n928);
   U5542 : AO6 port map( A => n930, B => n4789, C => n931, Z => n929);
   U5543 : AO3 port map( A => n4888, B => n4488, C => n107, D => n108, Z => 
                           n4071);
   U5544 : AO2 port map( A => n4785, B => n135, C => n136, D => n4787, Z => 
                           n107);
   U5545 : AO6 port map( A => n109, B => n4791, C => n111, Z => n108);
   U5546 : AO3 port map( A => n4887, B => n4489, C => n887, D => n888, Z => 
                           n4077);
   U5547 : AO2 port map( A => n4783, B => n917, C => n918, D => n4788, Z => 
                           n887);
   U5548 : AO6 port map( A => n889, B => n4789, C => n890, Z => n888);
   U5549 : AO3 port map( A => n4887, B => n4490, C => n423, D => n424, Z => 
                           n4084);
   U5550 : AO2 port map( A => n4784, B => n453, C => n454, D => n4787, Z => 
                           n423);
   U5551 : AO6 port map( A => n425, B => n4790, C => n426, Z => n424);
   U5552 : AO3 port map( A => n4886, B => n4493, C => n1065, D => n1066, Z => 
                           n4102);
   U5553 : AO2 port map( A => n4783, B => n1091, C => n1092, D => n4788, Z => 
                           n1065);
   U5554 : AO6 port map( A => n1067, B => n4789, C => n1068, Z => n1066);
   U5555 : AO3 port map( A => n4887, B => n4494, C => n725, D => n726, Z => 
                           n4108);
   U5556 : AO2 port map( A => n4783, B => n746, C => n747, D => n4788, Z => 
                           n725);
   U5557 : AO6 port map( A => n727, B => n4789, C => n728, Z => n726);
   U5558 : AO3 port map( A => n4888, B => n4495, C => n233, D => n234, Z => 
                           n4115);
   U5559 : AO2 port map( A => n4784, B => n257, C => n258, D => n4787, Z => 
                           n233);
   U5560 : AO6 port map( A => n235, B => n4790, C => n236, Z => n234);
   U5561 : AO3 port map( A => n4886, B => n4496, C => n1038, D => n1039, Z => 
                           n4121);
   U5562 : AO2 port map( A => n4783, B => n1058, C => n1059, D => n4788, Z => 
                           n1038);
   U5563 : AO6 port map( A => n1040, B => n4789, C => n1041, Z => n1039);
   U5564 : AO3 port map( A => n4887, B => n4497, C => n696, D => n697, Z => 
                           n4127);
   U5565 : AO2 port map( A => n4783, B => n717, C => n718, D => n4788, Z => 
                           n696);
   U5566 : AO6 port map( A => n698, B => n4789, C => n699, Z => n697);
   U5567 : AO3 port map( A => n4888, B => n4498, C => n394, D => n395, Z => 
                           n4133);
   U5568 : AO2 port map( A => n4784, B => n415, C => n416, D => n4787, Z => 
                           n394);
   U5569 : AO6 port map( A => n396, B => n4790, C => n397, Z => n395);
   U5570 : AO3 port map( A => n4888, B => n4499, C => n204, D => n205, Z => 
                           n4140);
   U5571 : AO2 port map( A => n4784, B => n225, C => n226, D => n4787, Z => 
                           n204);
   U5572 : AO6 port map( A => n206, B => n4790, C => n207, Z => n205);
   U5573 : AO3 port map( A => n4886, B => n4500, C => n1009, D => n1010, Z => 
                           n4146);
   U5574 : AO2 port map( A => n4783, B => n1031, C => n1032, D => n4788, Z => 
                           n1009);
   U5575 : AO6 port map( A => n1011, B => n4789, C => n1012, Z => n1010);
   U5576 : AO3 port map( A => n4887, B => n4501, C => n663, D => n664, Z => 
                           n4152);
   U5577 : AO2 port map( A => n4783, B => n687, C => n688, D => n4788, Z => 
                           n663);
   U5578 : AO6 port map( A => n665, B => n4789, C => n666, Z => n664);
   U5579 : AO3 port map( A => n4888, B => n4502, C => n373, D => n374, Z => 
                           n4158);
   U5580 : AO2 port map( A => n4784, B => n388, C => n389, D => n4787, Z => 
                           n373);
   U5581 : AO6 port map( A => n375, B => n4790, C => n376, Z => n374);
   U5582 : AO3 port map( A => n4887, B => n4503, C => n620, D => n621, Z => 
                           n4165);
   U5583 : AO2 port map( A => n4784, B => n651, C => n652, D => n4788, Z => 
                           n620);
   U5584 : AO6 port map( A => n622, B => n4790, C => n623, Z => n621);
   U5585 : NR3 port map( A => n5023, B => RESET_I, C => n1301, Z => n1315);
   U5586 : AO7 port map( A => n3827, B => n4743, C => n4952, Z => n4174);
   U5587 : AO4 port map( A => n1967, B => n5065, C => n4840, D => n296, Z => 
                           n1976);
   U5588 : AO7 port map( A => n3828, B => n4744, C => n4950, Z => n4175);
   U5589 : AO4 port map( A => n1967, B => n1618, C => n4840, D => n261, Z => 
                           n1974);
   U5590 : AO7 port map( A => n3843, B => n4734, C => n4923, Z => n4190);
   U5591 : AO4 port map( A => n2410, B => n5073, C => n4842, D => n264, Z => 
                           n2419);
   U5592 : NR3 port map( A => n3954, B => n5005, C => n5011, Z => n1430);
   U5593 : AO4 port map( A => n3958, B => n5020, C => n4439, D => n1444, Z => 
                           n1418);
   U5594 : AO7 port map( A => n3957, B => n1418, C => CE_I, Z => n1441);
   U5595 : AO3 port map( A => n1601, B => n1893, C => n1935, D => n1936, Z => 
                           n4078);
   U5596 : AO3 port map( A => n1595, B => n1893, C => n1912, D => n1913, Z => 
                           n4109);
   U5597 : AO3 port map( A => n1584, B => n1893, C => n1905, D => n1906, Z => 
                           n4159);
   U5598 : AO3 port map( A => n1557, B => n2410, C => n2452, D => n2453, Z => 
                           n4186);
   U5599 : AO3 port map( A => n1545, B => n2410, C => n2424, D => n2425, Z => 
                           n4188);
   U5600 : AO3 port map( A => n1539, B => n2410, C => n2420, D => n2421, Z => 
                           n4189);
   U5601 : AO3 port map( A => n1805, B => n2888, C => n3186, D => n3187, Z => 
                           n4203);
   U5602 : AO3 port map( A => n1632, B => n2888, C => n3142, D => n3143, Z => 
                           n4204);
   U5603 : AO7 port map( A => n3956, B => n1428, C => n1429, Z => n4289);
   U5604 : AO6 port map( A => n3955, B => n1433, C => n1434, Z => n1428);
   U5605 : ND4 port map( A => n3956, B => n1430, C => n4633, D => n4471, Z => 
                           n1429);
   U5606 : EON1 port map( A => n3953, B => n1436, C => n1430, D => n3953, Z => 
                           n4291);
   U5607 : ND2I port map( A => v_RAM_OUT0_19_port, B => n4512, Z => n2982);
   U5608 : ND2I port map( A => v_RAM_OUT0_3_port, B => n4511, Z => n3385);
   U5609 : NR4 port map( A => n4411, B => v_CALCULATION_CNTR_3_port, C => n4527
                           , D => n3812, Z => n3805);
   U5610 : IVDA port map( A => v_RAM_OUT0_28_port, Y => n4360, Z => n4781);
   U5611 : IVDA port map( A => v_RAM_OUT0_20_port, Y => n4355, Z => n4780);
   U5612 : IVDA port map( A => v_RAM_OUT0_4_port, Y => n4358, Z => n4779);
   U5613 : AO3 port map( A => n1562, B => n1727, C => n1754, D => n1755, Z => 
                           n4249);
   U5614 : AO3 port map( A => n1557, B => n1727, C => n1750, D => n1751, Z => 
                           n4250);
   U5615 : AO3 port map( A => n1551, B => n1727, C => n1746, D => n1747, Z => 
                           n4251);
   U5616 : AO3 port map( A => n1545, B => n1727, C => n1742, D => n1743, Z => 
                           n4252);
   U5617 : AO3 port map( A => n1539, B => n1727, C => n1738, D => n1739, Z => 
                           n4253);
   U5618 : ND2I port map( A => v_RAM_OUT0_11_port, B => n4533, Z => n2033);
   U5619 : ND2I port map( A => v_RAM_OUT0_27_port, B => n4532, Z => n2575);
   U5620 : ND2I port map( A => v_RAM_OUT0_22_port, B => n4373, Z => n3015);
   U5621 : ND2I port map( A => v_RAM_OUT0_6_port, B => n4372, Z => n3418);
   U5622 : AO4 port map( A => n3902, B => n5017, C => n3910, D => n5019, Z => 
                           n3797);
   U5623 : AO7 port map( A => n3814, B => n5020, C => n3801, Z => n3796);
   U5624 : AO2 port map( A => n4701, B => n4573, C => n4702, D => n4462, Z => 
                           n3801);
   U5625 : AO4 port map( A => n3903, B => n5017, C => n3911, D => n5019, Z => 
                           n3786);
   U5626 : AO7 port map( A => n3815, B => n5020, C => n3787, Z => n3785);
   U5627 : AO2 port map( A => n4701, B => n4559, C => n4702, D => n4443, Z => 
                           n3787);
   U5628 : AO4 port map( A => n3904, B => n5017, C => n3912, D => n5019, Z => 
                           n3775);
   U5629 : AO7 port map( A => n3816, B => n5020, C => n3776, Z => n3774);
   U5630 : AO2 port map( A => n4701, B => n4574, C => n4702, D => n4436, Z => 
                           n3776);
   U5631 : AO4 port map( A => n3905, B => n5017, C => n3913, D => n5019, Z => 
                           n3764);
   U5632 : AO7 port map( A => n3817, B => n5020, C => n3765, Z => n3763);
   U5633 : AO2 port map( A => n4701, B => n4575, C => n4702, D => n4452, Z => 
                           n3765);
   U5634 : AO4 port map( A => n3906, B => n5017, C => n3914, D => n5019, Z => 
                           n3753);
   U5635 : AO7 port map( A => n3818, B => n5020, C => n3754, Z => n3752);
   U5636 : AO2 port map( A => n4701, B => n4560, C => n4702, D => n4453, Z => 
                           n3754);
   U5637 : AO4 port map( A => n3907, B => n5017, C => n3915, D => n5019, Z => 
                           n3742);
   U5638 : AO7 port map( A => n3819, B => n5020, C => n3743, Z => n3741);
   U5639 : AO2 port map( A => n4701, B => n4408, C => n4702, D => n4572, Z => 
                           n3743);
   U5640 : AO4 port map( A => n3908, B => n5017, C => n3916, D => n5019, Z => 
                           n3730);
   U5641 : AO7 port map( A => n3820, B => n5020, C => n3731, Z => n3729);
   U5642 : AO2 port map( A => n4701, B => n4437, C => n4702, D => n4384, Z => 
                           n3731);
   U5643 : AO4 port map( A => n3909, B => n5017, C => n3917, D => n5019, Z => 
                           n3717);
   U5644 : AO7 port map( A => n3821, B => n5020, C => n3720, Z => n3716);
   U5645 : AO2 port map( A => n4701, B => n4548, C => n4702, D => n4420, Z => 
                           n3720);
   U5646 : AO3 port map( A => n4365, B => n2200, C => v_RAM_OUT0_13_port, D => 
                           n2356, Z => n2352);
   U5647 : AO6 port map( A => n4515, B => v_RAM_OUT0_11_port, C => n2357, Z => 
                           n2356);
   U5648 : AO4 port map( A => n2059, B => n4376, C => n4737, D => n2358, Z => 
                           n2357);
   U5649 : AO3 port map( A => n1601, B => n1758, C => n1780, D => n1781, Z => 
                           n4258);
   U5650 : AO3 port map( A => n1595, B => n1758, C => n1776, D => n1777, Z => 
                           n4259);
   U5651 : AO3 port map( A => n1584, B => n1758, C => n1769, D => n1770, Z => 
                           n4261);
   U5652 : AO3 port map( A => n1787, B => n1813, C => n1814, D => n1815, Z => 
                           n4265);
   U5653 : AO3 port map( A => n1787, B => n1805, C => n1806, D => n1807, Z => 
                           n4267);
   U5654 : AO3 port map( A => n1632, B => n1787, C => n1801, D => n1802, Z => 
                           n4268);
   U5655 : AO4 port map( A => n3954, B => n1439, C => n5005, D => n1440, Z => 
                           n4292);
   U5656 : EON1 port map( A => n4527, B => n1413, C => N2086, D => n1409, Z => 
                           n4309);
   U5657 : EON1 port map( A => n4556, B => n1413, C => N2084, D => n1409, Z => 
                           n4311);
   U5658 : EOI port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => N2083);
   U5659 : EON1 port map( A => n4604, B => n1413, C => n4604, D => n1409, Z => 
                           n4313);
   U5660 : AO3 port map( A => n3918, B => n4841, C => n3789, D => n3790, Z => 
                           n3961);
   U5661 : AO2 port map( A => n4854, B => n4610, C => n4692, D => DATA_O_0_port
                           , Z => n3790);
   U5662 : AO2 port map( A => n4353, B => n3791, C => n4848, D => n4605, Z => 
                           n3789);
   U5663 : ND4 port map( A => n3792, B => n3793, C => n3794, D => n3795, Z => 
                           n3791);
   U5664 : AO3 port map( A => n3919, B => n4841, C => n3778, D => n3779, Z => 
                           n3962);
   U5665 : AO2 port map( A => n4854, B => n4611, C => n4692, D => DATA_O_1_port
                           , Z => n3779);
   U5666 : AO2 port map( A => n4352, B => n3780, C => n4848, D => n4606, Z => 
                           n3778);
   U5667 : ND4 port map( A => n3781, B => n3782, C => n3783, D => n3784, Z => 
                           n3780);
   U5668 : AO3 port map( A => n3920, B => n4842, C => n3767, D => n3768, Z => 
                           n3963);
   U5669 : AO2 port map( A => n4854, B => n4418, C => n4692, D => DATA_O_2_port
                           , Z => n3768);
   U5670 : AO2 port map( A => n4353, B => n3769, C => n4848, D => n4607, Z => 
                           n3767);
   U5671 : ND4 port map( A => n3770, B => n3771, C => n3772, D => n3773, Z => 
                           n3769);
   U5672 : AO3 port map( A => n3921, B => n4842, C => n3756, D => n3757, Z => 
                           n3964);
   U5673 : AO2 port map( A => n4854, B => n4442, C => n4692, D => DATA_O_3_port
                           , Z => n3757);
   U5674 : AO2 port map( A => n4352, B => n3758, C => n4848, D => n4608, Z => 
                           n3756);
   U5675 : ND4 port map( A => n3759, B => n3760, C => n3761, D => n3762, Z => 
                           n3758);
   U5676 : AO3 port map( A => n3922, B => n4842, C => n3745, D => n3746, Z => 
                           n3965);
   U5677 : AO2 port map( A => n4854, B => n4551, C => n4692, D => DATA_O_4_port
                           , Z => n3746);
   U5678 : AO2 port map( A => n4353, B => n3747, C => n4848, D => n4609, Z => 
                           n3745);
   U5679 : ND4 port map( A => n3748, B => n3749, C => n3750, D => n3751, Z => 
                           n3747);
   U5680 : AO3 port map( A => n3923, B => n4842, C => n3734, D => n3735, Z => 
                           n3966);
   U5681 : AO2 port map( A => n4854, B => n4612, C => n4691, D => DATA_O_5_port
                           , Z => n3735);
   U5682 : AO2 port map( A => n4352, B => n3736, C => n4848, D => n4523, Z => 
                           n3734);
   U5683 : ND4 port map( A => n3737, B => n3738, C => n3739, D => n3740, Z => 
                           n3736);
   U5684 : AO3 port map( A => n3924, B => n4842, C => n3722, D => n3723, Z => 
                           n3967);
   U5685 : AO2 port map( A => n4854, B => n4419, C => n4691, D => DATA_O_6_port
                           , Z => n3723);
   U5686 : AO2 port map( A => n4353, B => n3724, C => n4848, D => n4406, Z => 
                           n3722);
   U5687 : ND4 port map( A => n3725, B => n3726, C => n3727, D => n3728, Z => 
                           n3724);
   U5688 : AO3 port map( A => n3925, B => n4841, C => n3705, D => n3706, Z => 
                           n3968);
   U5689 : AO2 port map( A => n4854, B => n4407, C => n4691, D => DATA_O_7_port
                           , Z => n3706);
   U5690 : AO2 port map( A => n4352, B => n3710, C => n4848, D => n4431, Z => 
                           n3705);
   U5691 : ND4 port map( A => n3712, B => n3713, C => n3714, D => n3715, Z => 
                           n3710);
   U5692 : AO2 port map( A => n5009, B => v_CALCULATION_CNTR_7_port, C => N2089
                           , D => n1409, Z => n1407);
   U5693 : AO2 port map( A => n5009, B => v_CALCULATION_CNTR_6_port, C => N2088
                           , D => n1409, Z => n1410);
   U5694 : AO2 port map( A => n5009, B => v_CALCULATION_CNTR_5_port, C => N2087
                           , D => n1409, Z => n1411);
   U5695 : NR4 port map( A => n2377, B => n4527, C => n3809, D => 
                           v_CALCULATION_CNTR_5_port, Z => n3804);
   U5696 : AO6 port map( A => v_RAM_OUT0_11_port, B => n4552, C => n2078, Z => 
                           n2272);
   U5697 : AO4 port map( A => n3813, B => n4855, C => n3958, D => n1460, Z => 
                           n3960);
   U5698 : NR4 port map( A => n4701, B => n4700, C => n1478, D => n1479, Z => 
                           n1461);
   U5699 : NR4 port map( A => n5021, B => n1353, C => n1474, D => n4702, Z => 
                           n1462);
   U5700 : ND2I port map( A => v_RAM_OUT0_30_port, B => n4374, Z => n2609);
   U5701 : IVDA port map( A => v_RAM_OUT0_21_port, Y => n4403, Z => n4782);
   U5702 : AO6 port map( A => n4697, B => n4547, C => n3803, Z => n3794);
   U5703 : AO4 port map( A => n3838, B => n4698, C => n3854, D => n4699, Z => 
                           n3803);
   U5704 : AO6 port map( A => n4697, B => n4586, C => n3788, Z => n3783);
   U5705 : AO4 port map( A => n3839, B => n4698, C => n3855, D => n4699, Z => 
                           n3788);
   U5706 : AO6 port map( A => n4697, B => n4587, C => n3777, Z => n3772);
   U5707 : AO4 port map( A => n3840, B => n4698, C => n3856, D => n4699, Z => 
                           n3777);
   U5708 : AO6 port map( A => n4697, B => n4588, C => n3766, Z => n3761);
   U5709 : AO4 port map( A => n3841, B => n4698, C => n3857, D => n4699, Z => 
                           n3766);
   U5710 : AO6 port map( A => n4697, B => n4558, C => n3755, Z => n3750);
   U5711 : AO4 port map( A => n3842, B => n4698, C => n3858, D => n4699, Z => 
                           n3755);
   U5712 : AO6 port map( A => n4697, B => n4541, C => n3744, Z => n3739);
   U5713 : AO4 port map( A => n3843, B => n4698, C => n3859, D => n4699, Z => 
                           n3744);
   U5714 : AO6 port map( A => n4697, B => n4598, C => n3733, Z => n3727);
   U5715 : AO4 port map( A => n3844, B => n4698, C => n3860, D => n4699, Z => 
                           n3733);
   U5716 : AO6 port map( A => n4697, B => n4589, C => n3721, Z => n3714);
   U5717 : AO4 port map( A => n3845, B => n4698, C => n3861, D => n4699, Z => 
                           n3721);
   U5718 : AO3 port map( A => n3957, B => n1413, C => n3810, D => n3811, Z => 
                           n4293);
   U5719 : ND4 port map( A => CE_I, B => n5010, C => n4999, D => n4414, Z => 
                           n3811);
   U5720 : AO7 port map( A => n3958, B => n5020, C => n1433, Z => n3810);
   U5721 : AO7 port map( A => n1433, B => n5009, C => n4439, Z => n3700);
   U5722 : ND4 port map( A => n3953, B => n5022, C => n5012, D => n3703, Z => 
                           n3701);
   U5723 : NR3 port map( A => n3956, B => n3955, C => n4892, Z => n3703);
   U5724 : AO3 port map( A => n4764, B => n3947, C => n1355, D => n1356, Z => 
                           n4301);
   U5725 : EON1 port map( A => n4472, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_0_port, Z => n3972);
   U5726 : EON1 port map( A => n4473, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_16_port, Z => n3978);
   U5727 : EON1 port map( A => n4474, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_8_port, Z => n3984);
   U5728 : EON1 port map( A => n4475, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_3_port, Z => n3990);
   U5729 : EON1 port map( A => n4476, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_11_port, Z => n3996);
   U5730 : EON1 port map( A => n4477, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_19_port, Z => n4002);
   U5731 : EON1 port map( A => n4478, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_27_port, Z => n4008);
   U5732 : EON1 port map( A => n4479, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_10_port, Z => n4014);
   U5733 : EON1 port map( A => n4480, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_26_port, Z => n4020);
   U5734 : EON1 port map( A => n4481, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_17_port, Z => n4026);
   U5735 : EON1 port map( A => n4482, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_25_port, Z => n4032);
   U5736 : EON1 port map( A => n4483, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_1_port, Z => n4039);
   U5737 : EON1 port map( A => n4484, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_4_port, Z => n4045);
   U5738 : EON1 port map( A => n4485, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_20_port, Z => n4051);
   U5739 : EON1 port map( A => n4486, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_12_port, Z => n4057);
   U5740 : EON1 port map( A => n4487, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_28_port, Z => n4063);
   U5741 : EON1 port map( A => n4488, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_9_port, Z => n4069);
   U5742 : EON1 port map( A => n4489, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_18_port, Z => n4075);
   U5743 : EON1 port map( A => n4490, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_2_port, Z => n4082);
   U5744 : EON1 port map( A => n4491, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_5_port, Z => n4088);
   U5745 : EON1 port map( A => n4492, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_29_port, Z => n4094);
   U5746 : EON1 port map( A => n4493, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_13_port, Z => n4100);
   U5747 : EON1 port map( A => n4494, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_21_port, Z => n4106);
   U5748 : EON1 port map( A => n4495, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_6_port, Z => n4113);
   U5749 : EON1 port map( A => n4496, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_14_port, Z => n4119);
   U5750 : EON1 port map( A => n4497, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_22_port, Z => n4125);
   U5751 : EON1 port map( A => n4498, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_30_port, Z => n4131);
   U5752 : EON1 port map( A => n4499, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_7_port, Z => n4138);
   U5753 : EON1 port map( A => n4500, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_15_port, Z => n4144);
   U5754 : EON1 port map( A => n4501, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_23_port, Z => n4150);
   U5755 : EON1 port map( A => n4502, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_31_port, Z => n4156);
   U5756 : EON1 port map( A => n4503, B => n4361, C => n4361, D => 
                           t_STATE_RAM0_1_24_port, Z => n4163);
   U5757 : IVDA port map( A => n1354, Y => n_3431, Z => n4764);
   U5758 : AO7 port map( A => n3952, B => n4892, C => n5002, Z => n1354);
   U5759 : AO7 port map( A => n4764, B => n3946, C => n1359, Z => n4298);
   U5760 : ND4 port map( A => N200, B => n4764, C => n1360, D => n5010, Z => 
                           n1359);
   U5761 : AO7 port map( A => n5000, B => RESET_I, C => n4764, Z => n1355);
   U5762 : ND4 port map( A => CE_I, B => n1458, C => n4556, D => n4369, Z => 
                           n1452);
   U5763 : AO3 port map( A => n4764, B => n3944, C => n1355, D => n1357, Z => 
                           n4296);
   U5764 : AO3 port map( A => n4367, B => n4634, C => n100, D => n101, Z => 
                           n3969);
   U5765 : AO2 port map( A => t_STATE_RAM0_0_0_port, B => n4891, C => 
                           t_STATE_RAM0_2_0_port, D => n4890, Z => n100);
   U5766 : AO2 port map( A => t_STATE_RAM0_1_0_port, B => n4363, C => 
                           v_RAM_OUT0_0_port, D => n4892, Z => n101);
   U5767 : EON1 port map( A => n4472, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_0_port, Z => n3971);
   U5768 : EON1 port map( A => n4472, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_0_port, Z => n3973);
   U5769 : AO3 port map( A => n4367, B => n4635, C => n79, D => n80, Z => n3975
                           );
   U5770 : AO2 port map( A => t_STATE_RAM0_0_16_port, B => n4891, C => 
                           t_STATE_RAM0_2_16_port, D => n4890, Z => n79);
   U5771 : AO2 port map( A => t_STATE_RAM0_1_16_port, B => n4363, C => 
                           v_RAM_OUT0_16_port, D => n4892, Z => n80);
   U5772 : EON1 port map( A => n4473, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_16_port, Z => n3977);
   U5773 : EON1 port map( A => n4473, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_16_port, Z => n3979);
   U5774 : AO3 port map( A => n4367, B => n4636, C => n10, D => n11, Z => n3981
                           );
   U5775 : AO2 port map( A => t_STATE_RAM0_0_8_port, B => n4891, C => 
                           t_STATE_RAM0_2_8_port, D => n4890, Z => n10);
   U5776 : AO2 port map( A => t_STATE_RAM0_1_8_port, B => n4363, C => n4775, D 
                           => n4892, Z => n11);
   U5777 : EON1 port map( A => n4474, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_8_port, Z => n3983);
   U5778 : EON1 port map( A => n4474, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_8_port, Z => n3985);
   U5779 : AO3 port map( A => n4367, B => n4637, C => n25, D => n26, Z => n3987
                           );
   U5780 : AO2 port map( A => t_STATE_RAM0_0_3_port, B => n4891, C => 
                           t_STATE_RAM0_2_3_port, D => n4890, Z => n25);
   U5781 : AO2 port map( A => t_STATE_RAM0_1_3_port, B => n4363, C => 
                           v_RAM_OUT0_3_port, D => n4892, Z => n26);
   U5782 : EON1 port map( A => n4475, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_3_port, Z => n3989);
   U5783 : EON1 port map( A => n4475, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_3_port, Z => n3991);
   U5784 : AO3 port map( A => n4367, B => n4638, C => n94, D => n95, Z => n3993
                           );
   U5785 : AO2 port map( A => t_STATE_RAM0_0_11_port, B => n4891, C => 
                           t_STATE_RAM0_2_11_port, D => n4890, Z => n94);
   U5786 : AO2 port map( A => t_STATE_RAM0_1_11_port, B => n4363, C => 
                           v_RAM_OUT0_11_port, D => n4892, Z => n95);
   U5787 : EON1 port map( A => n4476, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_11_port, Z => n3995);
   U5788 : EON1 port map( A => n4476, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_11_port, Z => n3997);
   U5789 : AO3 port map( A => n4367, B => n4639, C => n70, D => n71, Z => n3999
                           );
   U5790 : AO2 port map( A => t_STATE_RAM0_0_19_port, B => n4891, C => 
                           t_STATE_RAM0_2_19_port, D => n4890, Z => n70);
   U5791 : AO2 port map( A => t_STATE_RAM0_1_19_port, B => n4363, C => 
                           v_RAM_OUT0_19_port, D => n4892, Z => n71);
   U5792 : EON1 port map( A => n4477, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_19_port, Z => n4001);
   U5793 : EON1 port map( A => n4477, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_19_port, Z => n4003);
   U5794 : AO3 port map( A => n4367, B => n4640, C => n43, D => n44, Z => n4005
                           );
   U5795 : AO2 port map( A => t_STATE_RAM0_0_27_port, B => n4891, C => 
                           t_STATE_RAM0_2_27_port, D => n4890, Z => n43);
   U5796 : AO2 port map( A => t_STATE_RAM0_1_27_port, B => n4363, C => 
                           v_RAM_OUT0_27_port, D => n4892, Z => n44);
   U5797 : EON1 port map( A => n4478, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_27_port, Z => n4007);
   U5798 : EON1 port map( A => n4478, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_27_port, Z => n4009);
   U5799 : AO3 port map( A => n4367, B => n4641, C => n97, D => n98, Z => n4011
                           );
   U5800 : AO2 port map( A => t_STATE_RAM0_0_10_port, B => n4891, C => 
                           t_STATE_RAM0_2_10_port, D => n4890, Z => n97);
   U5801 : AO2 port map( A => t_STATE_RAM0_1_10_port, B => n4363, C => 
                           v_RAM_OUT0_10_port, D => n4892, Z => n98);
   U5802 : EON1 port map( A => n4479, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_10_port, Z => n4013);
   U5803 : EON1 port map( A => n4479, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_10_port, Z => n4015);
   U5804 : AO3 port map( A => n4367, B => n4642, C => n46, D => n47, Z => n4017
                           );
   U5805 : AO2 port map( A => t_STATE_RAM0_0_26_port, B => n4891, C => 
                           t_STATE_RAM0_2_26_port, D => n4890, Z => n46);
   U5806 : AO2 port map( A => t_STATE_RAM0_1_26_port, B => n4363, C => 
                           v_RAM_OUT0_26_port, D => n4892, Z => n47);
   U5807 : EON1 port map( A => n4480, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_26_port, Z => n4019);
   U5808 : EON1 port map( A => n4480, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_26_port, Z => n4021);
   U5809 : AO3 port map( A => n4367, B => n4643, C => n76, D => n77, Z => n4023
                           );
   U5810 : AO2 port map( A => t_STATE_RAM0_0_17_port, B => n4891, C => 
                           t_STATE_RAM0_2_17_port, D => n4890, Z => n76);
   U5811 : AO2 port map( A => t_STATE_RAM0_1_17_port, B => n4363, C => 
                           v_RAM_OUT0_17_port, D => n4892, Z => n77);
   U5812 : EON1 port map( A => n4481, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_17_port, Z => n4025);
   U5813 : EON1 port map( A => n4481, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_17_port, Z => n4027);
   U5814 : AO3 port map( A => n4367, B => n4644, C => n49, D => n50, Z => n4029
                           );
   U5815 : AO2 port map( A => t_STATE_RAM0_0_25_port, B => n4891, C => 
                           t_STATE_RAM0_2_25_port, D => n4890, Z => n49);
   U5816 : AO2 port map( A => t_STATE_RAM0_1_25_port, B => n4363, C => 
                           v_RAM_OUT0_25_port, D => n4892, Z => n50);
   U5817 : EON1 port map( A => n4482, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_25_port, Z => n4031);
   U5818 : EON1 port map( A => n4482, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_25_port, Z => n4033);
   U5819 : AO3 port map( A => n4367, B => n4645, C => n67, D => n68, Z => n4036
                           );
   U5820 : AO2 port map( A => t_STATE_RAM0_0_1_port, B => n4891, C => 
                           t_STATE_RAM0_2_1_port, D => n4890, Z => n67);
   U5821 : AO2 port map( A => t_STATE_RAM0_1_1_port, B => n4363, C => 
                           v_RAM_OUT0_1_port, D => n4892, Z => n68);
   U5822 : EON1 port map( A => n4483, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_1_port, Z => n4038);
   U5823 : EON1 port map( A => n4483, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_1_port, Z => n4040);
   U5824 : AO3 port map( A => n4367, B => n4646, C => n22, D => n23, Z => n4042
                           );
   U5825 : AO2 port map( A => t_STATE_RAM0_0_4_port, B => n4891, C => 
                           t_STATE_RAM0_2_4_port, D => n4890, Z => n22);
   U5826 : AO2 port map( A => t_STATE_RAM0_1_4_port, B => n4363, C => n4779, D 
                           => n4892, Z => n23);
   U5827 : EON1 port map( A => n4484, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_4_port, Z => n4044);
   U5828 : EON1 port map( A => n4484, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_4_port, Z => n4046);
   U5829 : AO3 port map( A => n4367, B => n4647, C => n64, D => n65, Z => n4048
                           );
   U5830 : AO2 port map( A => t_STATE_RAM0_0_20_port, B => n4891, C => 
                           t_STATE_RAM0_2_20_port, D => n4890, Z => n64);
   U5831 : AO2 port map( A => t_STATE_RAM0_1_20_port, B => n4363, C => n4780, D
                           => n4892, Z => n65);
   U5832 : EON1 port map( A => n4485, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_20_port, Z => n4050);
   U5833 : EON1 port map( A => n4485, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_20_port, Z => n4052);
   U5834 : AO3 port map( A => n4367, B => n4648, C => n91, D => n92, Z => n4054
                           );
   U5835 : AO2 port map( A => t_STATE_RAM0_0_12_port, B => n4891, C => 
                           t_STATE_RAM0_2_12_port, D => n4890, Z => n91);
   U5836 : AO2 port map( A => t_STATE_RAM0_1_12_port, B => n4363, C => 
                           v_RAM_OUT0_12_port, D => n4892, Z => n92);
   U5837 : EON1 port map( A => n4486, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_12_port, Z => n4056);
   U5838 : EON1 port map( A => n4486, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_12_port, Z => n4058);
   U5839 : AO3 port map( A => n4367, B => n4649, C => n40, D => n41, Z => n4060
                           );
   U5840 : AO2 port map( A => t_STATE_RAM0_0_28_port, B => n4891, C => 
                           t_STATE_RAM0_2_28_port, D => n4890, Z => n40);
   U5841 : AO2 port map( A => t_STATE_RAM0_1_28_port, B => n4363, C => n4781, D
                           => n4892, Z => n41);
   U5842 : EON1 port map( A => n4487, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_28_port, Z => n4062);
   U5843 : EON1 port map( A => n4487, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_28_port, Z => n4064);
   U5844 : AO3 port map( A => n4367, B => n4650, C => n3, D => n4, Z => n4066);
   U5845 : AO2 port map( A => t_STATE_RAM0_0_9_port, B => n4891, C => 
                           t_STATE_RAM0_2_9_port, D => n4890, Z => n3);
   U5846 : AO2 port map( A => t_STATE_RAM0_1_9_port, B => n4363, C => 
                           v_RAM_OUT0_9_port, D => n4892, Z => n4);
   U5847 : EON1 port map( A => n4488, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_9_port, Z => n4068);
   U5848 : EON1 port map( A => n4488, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_9_port, Z => n4070);
   U5849 : AO3 port map( A => n4367, B => n4651, C => n73, D => n74, Z => n4072
                           );
   U5850 : AO2 port map( A => t_STATE_RAM0_0_18_port, B => n4891, C => 
                           t_STATE_RAM0_2_18_port, D => n4890, Z => n73);
   U5851 : AO2 port map( A => t_STATE_RAM0_1_18_port, B => n4363, C => 
                           v_RAM_OUT0_18_port, D => n4892, Z => n74);
   U5852 : EON1 port map( A => n4489, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_18_port, Z => n4074);
   U5853 : EON1 port map( A => n4489, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_18_port, Z => n4076);
   U5854 : AO3 port map( A => n4367, B => n4652, C => n34, D => n35, Z => n4079
                           );
   U5855 : AO2 port map( A => t_STATE_RAM0_0_2_port, B => n4891, C => 
                           t_STATE_RAM0_2_2_port, D => n4890, Z => n34);
   U5856 : AO2 port map( A => t_STATE_RAM0_1_2_port, B => n4363, C => 
                           v_RAM_OUT0_2_port, D => n4892, Z => n35);
   U5857 : EON1 port map( A => n4490, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_2_port, Z => n4081);
   U5858 : EON1 port map( A => n4490, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_2_port, Z => n4083);
   U5859 : AO3 port map( A => n4367, B => n4653, C => n19, D => n20, Z => n4085
                           );
   U5860 : AO2 port map( A => t_STATE_RAM0_0_5_port, B => n4891, C => 
                           t_STATE_RAM0_2_5_port, D => n4890, Z => n19);
   U5861 : AO2 port map( A => t_STATE_RAM0_1_5_port, B => n4363, C => 
                           v_RAM_OUT0_5_port, D => n4892, Z => n20);
   U5862 : EON1 port map( A => n4491, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_5_port, Z => n4087);
   U5863 : EON1 port map( A => n4491, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_5_port, Z => n4089);
   U5864 : AO3 port map( A => n4367, B => n4654, C => n37, D => n38, Z => n4091
                           );
   U5865 : AO2 port map( A => t_STATE_RAM0_0_29_port, B => n4891, C => 
                           t_STATE_RAM0_2_29_port, D => n4890, Z => n37);
   U5866 : AO2 port map( A => t_STATE_RAM0_1_29_port, B => n4363, C => 
                           v_RAM_OUT0_29_port, D => n4892, Z => n38);
   U5867 : EON1 port map( A => n4492, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_29_port, Z => n4093);
   U5868 : EON1 port map( A => n4492, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_29_port, Z => n4095);
   U5869 : AO3 port map( A => n4367, B => n4655, C => n88, D => n89, Z => n4097
                           );
   U5870 : AO2 port map( A => t_STATE_RAM0_0_13_port, B => n4891, C => 
                           t_STATE_RAM0_2_13_port, D => n4890, Z => n88);
   U5871 : AO2 port map( A => t_STATE_RAM0_1_13_port, B => n4363, C => 
                           v_RAM_OUT0_13_port, D => n4892, Z => n89);
   U5872 : EON1 port map( A => n4493, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_13_port, Z => n4099);
   U5873 : EON1 port map( A => n4493, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_13_port, Z => n4101);
   U5874 : AO3 port map( A => n4367, B => n4656, C => n61, D => n62, Z => n4103
                           );
   U5875 : AO2 port map( A => t_STATE_RAM0_0_21_port, B => n4891, C => 
                           t_STATE_RAM0_2_21_port, D => n4890, Z => n61);
   U5876 : AO2 port map( A => t_STATE_RAM0_1_21_port, B => n4363, C => n4782, D
                           => n4892, Z => n62);
   U5877 : EON1 port map( A => n4494, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_21_port, Z => n4105);
   U5878 : EON1 port map( A => n4494, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_21_port, Z => n4107);
   U5879 : AO3 port map( A => n4367, B => n4657, C => n16, D => n17, Z => n4110
                           );
   U5880 : AO2 port map( A => t_STATE_RAM0_0_6_port, B => n4891, C => 
                           t_STATE_RAM0_2_6_port, D => n4890, Z => n16);
   U5881 : AO2 port map( A => t_STATE_RAM0_1_6_port, B => n4363, C => 
                           v_RAM_OUT0_6_port, D => n4892, Z => n17);
   U5882 : EON1 port map( A => n4495, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_6_port, Z => n4112);
   U5883 : EON1 port map( A => n4495, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_6_port, Z => n4114);
   U5884 : AO3 port map( A => n4367, B => n4658, C => n85, D => n86, Z => n4116
                           );
   U5885 : AO2 port map( A => t_STATE_RAM0_0_14_port, B => n4891, C => 
                           t_STATE_RAM0_2_14_port, D => n4890, Z => n85);
   U5886 : AO2 port map( A => t_STATE_RAM0_1_14_port, B => n4363, C => 
                           v_RAM_OUT0_14_port, D => n4892, Z => n86);
   U5887 : EON1 port map( A => n4496, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_14_port, Z => n4118);
   U5888 : EON1 port map( A => n4496, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_14_port, Z => n4120);
   U5889 : AO3 port map( A => n4367, B => n4659, C => n58, D => n59, Z => n4122
                           );
   U5890 : AO2 port map( A => t_STATE_RAM0_0_22_port, B => n4891, C => 
                           t_STATE_RAM0_2_22_port, D => n4890, Z => n58);
   U5891 : AO2 port map( A => t_STATE_RAM0_1_22_port, B => n4363, C => 
                           v_RAM_OUT0_22_port, D => n4892, Z => n59);
   U5892 : EON1 port map( A => n4497, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_22_port, Z => n4124);
   U5893 : EON1 port map( A => n4497, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_22_port, Z => n4126);
   U5894 : AO3 port map( A => n4367, B => n4660, C => n31, D => n32, Z => n4128
                           );
   U5895 : AO2 port map( A => t_STATE_RAM0_0_30_port, B => n4891, C => 
                           t_STATE_RAM0_2_30_port, D => n4890, Z => n31);
   U5896 : AO2 port map( A => t_STATE_RAM0_1_30_port, B => n4363, C => 
                           v_RAM_OUT0_30_port, D => n4892, Z => n32);
   U5897 : EON1 port map( A => n4498, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_30_port, Z => n4130);
   U5898 : EON1 port map( A => n4498, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_30_port, Z => n4132);
   U5899 : AO3 port map( A => n4367, B => n4661, C => n13, D => n14, Z => n4135
                           );
   U5900 : AO2 port map( A => t_STATE_RAM0_0_7_port, B => n4891, C => 
                           t_STATE_RAM0_2_7_port, D => n4890, Z => n13);
   U5901 : AO2 port map( A => t_STATE_RAM0_1_7_port, B => n4363, C => 
                           v_RAM_OUT0_7_port, D => n4892, Z => n14);
   U5902 : EON1 port map( A => n4499, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_7_port, Z => n4137);
   U5903 : EON1 port map( A => n4499, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_7_port, Z => n4139);
   U5904 : AO3 port map( A => n4367, B => n4662, C => n82, D => n83, Z => n4141
                           );
   U5905 : AO2 port map( A => t_STATE_RAM0_0_15_port, B => n4891, C => 
                           t_STATE_RAM0_2_15_port, D => n4890, Z => n82);
   U5906 : AO2 port map( A => t_STATE_RAM0_1_15_port, B => n4363, C => 
                           v_RAM_OUT0_15_port, D => n4892, Z => n83);
   U5907 : EON1 port map( A => n4500, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_15_port, Z => n4143);
   U5908 : EON1 port map( A => n4500, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_15_port, Z => n4145);
   U5909 : AO3 port map( A => n4367, B => n4663, C => n55, D => n56, Z => n4147
                           );
   U5910 : AO2 port map( A => t_STATE_RAM0_0_23_port, B => n4891, C => 
                           t_STATE_RAM0_2_23_port, D => n4890, Z => n55);
   U5911 : AO2 port map( A => t_STATE_RAM0_1_23_port, B => n4363, C => 
                           v_RAM_OUT0_23_port, D => n4892, Z => n56);
   U5912 : EON1 port map( A => n4501, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_23_port, Z => n4149);
   U5913 : EON1 port map( A => n4501, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_23_port, Z => n4151);
   U5914 : AO3 port map( A => n4367, B => n4664, C => n28, D => n29, Z => n4153
                           );
   U5915 : AO2 port map( A => t_STATE_RAM0_0_31_port, B => n4891, C => 
                           t_STATE_RAM0_2_31_port, D => n4890, Z => n28);
   U5916 : AO2 port map( A => t_STATE_RAM0_1_31_port, B => n4363, C => 
                           v_RAM_OUT0_31_port, D => n4892, Z => n29);
   U5917 : EON1 port map( A => n4502, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_31_port, Z => n4155);
   U5918 : EON1 port map( A => n4502, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_31_port, Z => n4157);
   U5919 : AO3 port map( A => n4367, B => n4665, C => n52, D => n53, Z => n4160
                           );
   U5920 : AO2 port map( A => t_STATE_RAM0_0_24_port, B => n4891, C => 
                           t_STATE_RAM0_2_24_port, D => n4890, Z => n52);
   U5921 : AO2 port map( A => t_STATE_RAM0_1_24_port, B => n4363, C => 
                           v_RAM_OUT0_24_port, D => n4892, Z => n53);
   U5922 : EON1 port map( A => n4503, B => n4858, C => n4858, D => 
                           t_STATE_RAM0_2_24_port, Z => n4162);
   U5923 : EON1 port map( A => n4503, B => n4362, C => n4362, D => 
                           t_STATE_RAM0_0_24_port, Z => n4164);
   U5924 : AO3 port map( A => n4764, B => n3945, C => n1355, D => n1358, Z => 
                           n4297);
   U5925 : AO3 port map( A => n4666, B => n4764, C => n1355, D => n1361, Z => 
                           n4299);
   U5926 : AO3 port map( A => n4667, B => n4764, C => n1355, D => n1362, Z => 
                           n4300);
   U5927 : IVDA port map( A => n1377, Y => n4578, Z => n4763);
   U5928 : AO3 port map( A => CE_I, B => n4540, C => n1404, D => n4703, Z => 
                           n4340);
   U5929 : EON1 port map( A => n4998, B => n4763, C => n4763, D => 
                           v_DATA_COLUMN_24_port, Z => n4348);
   U5930 : IVDA port map( A => n1366, Y => n4465, Z => n4761);
   U5931 : AO2 port map( A => n4762, B => v_DATA_COLUMN_7_port, C => n4463, D 
                           => DATA_I(7), Z => n1369);
   U5932 : AO2 port map( A => n4762, B => v_DATA_COLUMN_6_port, C => n4463, D 
                           => DATA_I(6), Z => n1372);
   U5933 : AO2 port map( A => n4762, B => v_DATA_COLUMN_5_port, C => n4463, D 
                           => DATA_I(5), Z => n1373);
   U5934 : AO2 port map( A => n4762, B => v_DATA_COLUMN_4_port, C => n4463, D 
                           => DATA_I(4), Z => n1374);
   U5935 : AO2 port map( A => n4762, B => v_DATA_COLUMN_3_port, C => n4463, D 
                           => DATA_I(3), Z => n1375);
   U5936 : AO2 port map( A => n4762, B => v_DATA_COLUMN_2_port, C => n4463, D 
                           => DATA_I(2), Z => n1380);
   U5937 : AO2 port map( A => n4762, B => v_DATA_COLUMN_1_port, C => DATA_I(1),
                           D => n4463, Z => n1393);
   U5938 : AO2 port map( A => n4703, B => v_DATA_COLUMN_23_port, C => DATA_I(7)
                           , D => n4464, Z => n1387);
   U5939 : AO2 port map( A => n4703, B => v_DATA_COLUMN_22_port, C => DATA_I(6)
                           , D => n4464, Z => n1390);
   U5940 : AO2 port map( A => n4703, B => v_DATA_COLUMN_21_port, C => DATA_I(5)
                           , D => n4464, Z => n1391);
   U5941 : AO2 port map( A => n4703, B => v_DATA_COLUMN_20_port, C => DATA_I(4)
                           , D => n4464, Z => n1392);
   U5942 : AO2 port map( A => n4703, B => v_DATA_COLUMN_19_port, C => DATA_I(3)
                           , D => n4464, Z => n1394);
   U5943 : AO2 port map( A => n4703, B => v_DATA_COLUMN_18_port, C => DATA_I(2)
                           , D => n4464, Z => n1395);
   U5944 : AO2 port map( A => n4703, B => v_DATA_COLUMN_17_port, C => DATA_I(1)
                           , D => n4464, Z => n1396);
   U5945 : AO2 port map( A => n4761, B => v_DATA_COLUMN_15_port, C => n4465, D 
                           => DATA_I(7), Z => n1397);
   U5946 : AO2 port map( A => n4761, B => v_DATA_COLUMN_14_port, C => n4465, D 
                           => DATA_I(6), Z => n1398);
   U5947 : AO2 port map( A => n4761, B => v_DATA_COLUMN_13_port, C => n4465, D 
                           => DATA_I(5), Z => n1399);
   U5948 : AO2 port map( A => n4761, B => v_DATA_COLUMN_12_port, C => n4465, D 
                           => DATA_I(4), Z => n1400);
   U5949 : AO2 port map( A => n4761, B => v_DATA_COLUMN_11_port, C => n4465, D 
                           => DATA_I(3), Z => n1401);
   U5950 : AO2 port map( A => n4761, B => v_DATA_COLUMN_10_port, C => n4465, D 
                           => DATA_I(2), Z => n1402);
   U5951 : AO2 port map( A => n4761, B => v_DATA_COLUMN_9_port, C => n4465, D 
                           => DATA_I(1), Z => n1365);
   U5952 : AO2 port map( A => n4763, B => v_DATA_COLUMN_31_port, C => DATA_I(7)
                           , D => n4578, Z => n1376);
   U5953 : AO2 port map( A => n4763, B => v_DATA_COLUMN_30_port, C => DATA_I(6)
                           , D => n4578, Z => n1379);
   U5954 : AO2 port map( A => n4763, B => v_DATA_COLUMN_29_port, C => DATA_I(5)
                           , D => n4578, Z => n1381);
   U5955 : AO2 port map( A => n4763, B => v_DATA_COLUMN_28_port, C => DATA_I(4)
                           , D => n4578, Z => n1382);
   U5956 : AO2 port map( A => n4763, B => v_DATA_COLUMN_27_port, C => DATA_I(3)
                           , D => n4578, Z => n1383);
   U5957 : AO2 port map( A => n4763, B => v_DATA_COLUMN_26_port, C => n4578, D 
                           => DATA_I(2), Z => n1384);
   U5958 : AO2 port map( A => n4763, B => v_DATA_COLUMN_25_port, C => DATA_I(1)
                           , D => n4578, Z => n1385);
   U5959 : EON1 port map( A => n4999, B => n3704, C => n4414, D => n3704, Z => 
                           n4315);
   U5960 : AO4 port map( A => CE_I, B => n4380, C => n4999, D => n1406, Z => 
                           n4349);
   U5961 : AO4 port map( A => n3951, B => n4892, C => n3950, D => CE_I, Z => 
                           n4304);
   U5962 : AO4 port map( A => n3952, B => n4892, C => n3951, D => CE_I, Z => 
                           n4305);
   U5963 : IVI port map( A => CE_I, Z => n4892);
   U5964 : IVI port map( A => RESET_I, Z => n5010);
   U5965 : ND2I port map( A => n4779, B => n4371, Z => n4704);
   U5966 : ND2I port map( A => n4779, B => n4371, Z => n4705);
   U5967 : ND2I port map( A => v_RAM_OUT0_2_port, B => n4779, Z => n4707);
   U5968 : ND2I port map( A => v_RAM_OUT0_2_port, B => n4779, Z => n4708);
   U5969 : ND2I port map( A => n4780, B => n4395, Z => n4714);
   U5970 : ND2I port map( A => n4780, B => n4395, Z => n4715);
   U5971 : ND2I port map( A => v_RAM_OUT0_18_port, B => n4780, Z => n4717);
   U5972 : ND2I port map( A => v_RAM_OUT0_18_port, B => n4780, Z => n4718);
   U5973 : ND2I port map( A => v_RAM_OUT0_26_port, B => n4781, Z => n4725);
   U5974 : ND2I port map( A => v_RAM_OUT0_26_port, B => n4781, Z => n4726);
   U5975 : ND2I port map( A => n4781, B => n4397, Z => n4727);
   U5976 : ND2I port map( A => n4781, B => n4397, Z => n4728);
   U5977 : IVI port map( A => n4552, Z => n4771);
   U5978 : IVI port map( A => n4552, Z => n4772);
   U5979 : IVI port map( A => n4552, Z => n4773);
   U5980 : IVI port map( A => n4552, Z => n4774);
   U5981 : IVI port map( A => n4552, Z => n4775);
   U5982 : IVI port map( A => n4552, Z => n4776);
   U5983 : IVI port map( A => n4552, Z => n4777);
   U5984 : IVI port map( A => n4552, Z => n4778);
   U5985 : IVI port map( A => n4786, Z => n4785);
   U5986 : IVI port map( A => n5003, Z => n4786);
   U5987 : IVI port map( A => n4792, Z => n4791);
   U5988 : IVI port map( A => n5004, Z => n4792);
   U5989 : IVI port map( A => n4513, Z => n4793);
   U5990 : IVI port map( A => n4513, Z => n4794);
   U5991 : IVI port map( A => n4513, Z => n4795);
   U5992 : IVI port map( A => n4793, Z => n4798);
   U5993 : IVI port map( A => n4793, Z => n4799);
   U5994 : IVI port map( A => n4793, Z => n4800);
   U5995 : IVI port map( A => n4794, Z => n4801);
   U5996 : IVI port map( A => n4794, Z => n4802);
   U5997 : IVI port map( A => n4794, Z => n4803);
   U5998 : IVI port map( A => n4795, Z => n4804);
   U5999 : IVI port map( A => n4795, Z => n4805);
   U6000 : IVI port map( A => n3310, Z => n4808);
   U6001 : IVI port map( A => n4505, Z => n4809);
   U6002 : IVI port map( A => n4505, Z => n4810);
   U6003 : IVI port map( A => n4505, Z => n4811);
   U6004 : IVI port map( A => n4809, Z => n4814);
   U6005 : IVI port map( A => n4809, Z => n4815);
   U6006 : IVI port map( A => n4809, Z => n4816);
   U6007 : IVI port map( A => n4810, Z => n4817);
   U6008 : IVI port map( A => n4810, Z => n4818);
   U6009 : IVI port map( A => n4810, Z => n4819);
   U6010 : IVI port map( A => n4811, Z => n4820);
   U6011 : IVI port map( A => n4811, Z => n4821);
   U6012 : IVI port map( A => n4514, Z => n4824);
   U6013 : IVI port map( A => n4514, Z => n4825);
   U6014 : IVI port map( A => n4514, Z => n4826);
   U6015 : IVI port map( A => n4824, Z => n4829);
   U6016 : IVI port map( A => n4824, Z => n4830);
   U6017 : IVI port map( A => n4824, Z => n4831);
   U6018 : IVI port map( A => n4825, Z => n4832);
   U6019 : IVI port map( A => n4825, Z => n4833);
   U6020 : IVI port map( A => n4825, Z => n4834);
   U6021 : IVI port map( A => n4826, Z => n4835);
   U6022 : IVI port map( A => n4826, Z => n4836);
   U6023 : IVI port map( A => n1929, Z => n4839);
   U6024 : IVI port map( A => n4848, Z => n4847);
   U6025 : IVI port map( A => n1572, Z => n4848);
   U6026 : IVI port map( A => n4854, Z => n4853);
   U6027 : IVI port map( A => n1484, Z => n4854);
   U6028 : IVI port map( A => n4381, Z => n4857);
   U6029 : IVI port map( A => n4883, Z => n4859);
   U6030 : IVI port map( A => n4883, Z => n4860);
   U6031 : IVI port map( A => n4879, Z => n4861);
   U6032 : IVI port map( A => n4393, Z => n4862);
   U6033 : IVI port map( A => n4393, Z => n4863);
   U6034 : IVI port map( A => n4393, Z => n4864);
   U6035 : IVI port map( A => n4884, Z => n4867);
   U6036 : IVI port map( A => n4859, Z => n4868);
   U6037 : IVI port map( A => n4859, Z => n4869);
   U6038 : IVI port map( A => n4859, Z => n4870);
   U6039 : IVI port map( A => n4860, Z => n4871);
   U6040 : IVI port map( A => n4860, Z => n4872);
   U6041 : IVI port map( A => n4860, Z => n4873);
   U6042 : IVI port map( A => n4861, Z => n4874);
   U6043 : IVI port map( A => n4861, Z => n4875);
   U6044 : IVI port map( A => n4861, Z => n4876);
   U6045 : IVI port map( A => n4862, Z => n4877);
   U6046 : IVI port map( A => n4862, Z => n4878);
   U6047 : IVI port map( A => n4862, Z => n4879);
   U6048 : IVI port map( A => n4863, Z => n4880);
   U6049 : IVI port map( A => n4863, Z => n4881);
   U6050 : IVI port map( A => n4863, Z => n4882);
   U6051 : IVI port map( A => n4864, Z => n4883);
   U6052 : IVI port map( A => n4864, Z => n4884);
   U6053 : IVI port map( A => n105, Z => n4889);
   U6054 : IVI port map( A => n4584, Z => n4890);
   U6055 : IVI port map( A => n4585, Z => n4891);
   U6056 : ND2 port map( A => n4666, B => n4667, Z => n4893);
   U6057 : AO7 port map( A => n4667, B => n4666, C => n4893, Z => N199);
   U6058 : NR2 port map( A => n4893, B => v_INV_KEY_NUMB_2_port, Z => n4895);
   U6059 : AO6 port map( A => n4893, B => v_INV_KEY_NUMB_2_port, C => n4895, Z 
                           => n4894);
   U6060 : IV port map( A => n4894, Z => N200);
   U6061 : ND2 port map( A => n4895, B => n3945, Z => n4896);
   U6062 : AO7 port map( A => n4895, B => n3945, C => n4896, Z => N201);
   U6063 : EN port map( A => n4896, B => v_INV_KEY_NUMB_4_port, Z => N202);
   U6064 : NR2 port map( A => v_INV_KEY_NUMB_4_port, B => n4896, Z => n4897);
   U6065 : EO port map( A => v_INV_KEY_NUMB_5_port, B => n4897, Z => N203);
   U6066 : ND2 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n4898);
   U6067 : EN port map( A => n4898, B => v_CALCULATION_CNTR_2_port, Z => N2084)
                           ;
   U6068 : AN3 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, C => 
                           v_CALCULATION_CNTR_2_port, Z => n4900);
   U6069 : EO port map( A => n4900, B => v_CALCULATION_CNTR_3_port, Z => N2085)
                           ;
   U6070 : ND2 port map( A => v_CALCULATION_CNTR_3_port, B => n4900, Z => n4899
                           );
   U6071 : EN port map( A => n4899, B => v_CALCULATION_CNTR_4_port, Z => N2086)
                           ;
   U6072 : AN3 port map( A => v_CALCULATION_CNTR_3_port, B => n4900, C => 
                           v_CALCULATION_CNTR_4_port, Z => n4901);
   U6073 : EO port map( A => n4901, B => v_CALCULATION_CNTR_5_port, Z => N2087)
                           ;
   U6074 : ND2 port map( A => v_CALCULATION_CNTR_5_port, B => n4901, Z => n4902
                           );
   U6075 : EN port map( A => n4902, B => v_CALCULATION_CNTR_6_port, Z => N2088)
                           ;
   U6076 : NR2 port map( A => n4902, B => n4599, Z => n4903);
   U6077 : EO port map( A => v_CALCULATION_CNTR_7_port, B => n4903, Z => N2089)
                           ;
   U6078 : IVI port map( A => v_KEY_COLUMN_9_port, Z => n4904);
   U6079 : IVI port map( A => n449, Z => n4905);
   U6080 : IVI port map( A => n556, Z => n4906);
   U6081 : IVI port map( A => n831, Z => n4907);
   U6082 : IVI port map( A => n459, Z => n4908);
   U6083 : IVI port map( A => n546, Z => n4909);
   U6084 : IVI port map( A => n639, Z => n4910);
   U6085 : IVI port map( A => n999, Z => n4911);
   U6086 : IVI port map( A => n655, Z => n4912);
   U6087 : IVI port map( A => n630, Z => n4913);
   U6088 : IVI port map( A => n1088, Z => n4914);
   U6089 : IVI port map( A => n638, Z => n4915);
   U6090 : IVI port map( A => n1330, Z => n4916);
   U6091 : IVI port map( A => n1097, Z => n4917);
   U6092 : IVI port map( A => v_KEY_COLUMN_6_port, Z => n4918);
   U6093 : IVI port map( A => n1005, Z => n4919);
   U6094 : IVI port map( A => n1336, Z => n4920);
   U6095 : IVI port map( A => n231, Z => n4921);
   U6096 : IVI port map( A => v_KEY_COLUMN_5_port, Z => n4922);
   U6097 : IVI port map( A => n2419, Z => n4923);
   U6098 : IVI port map( A => n994, Z => n4924);
   U6099 : IVI port map( A => n612, Z => n4925);
   U6100 : IVI port map( A => n963, Z => n4926);
   U6101 : IVI port map( A => n1002, Z => n4927);
   U6102 : IVI port map( A => v_KEY_COLUMN_31_port, Z => n4928);
   U6103 : IVI port map( A => n673, Z => n4929);
   U6104 : IVI port map( A => n679, Z => n4930);
   U6105 : IVI port map( A => n685, Z => n4931);
   U6106 : IVI port map( A => n197, Z => n4932);
   U6107 : IVI port map( A => n968, Z => n4933);
   U6108 : IVI port map( A => n1019, Z => n4934);
   U6109 : IVI port map( A => n744, Z => n4935);
   U6110 : IVI port map( A => n1026, Z => n4936);
   U6111 : IVI port map( A => v_KEY_COLUMN_29_port, Z => n4937);
   U6112 : IVI port map( A => n780, Z => n4938);
   U6113 : IVI port map( A => n849, Z => n4939);
   U6114 : IVI port map( A => n860, Z => n4940);
   U6115 : IVI port map( A => n871, Z => n4941);
   U6116 : IVI port map( A => n884, Z => n4942);
   U6117 : IVI port map( A => n158, Z => n4943);
   U6118 : IVI port map( A => n183, Z => n4944);
   U6119 : IVI port map( A => n175, Z => n4945);
   U6120 : IVI port map( A => n192_port, Z => n4946);
   U6121 : IVI port map( A => n241, Z => n4947);
   U6122 : IVI port map( A => n253, Z => n4948);
   U6123 : IVI port map( A => n247, Z => n4949);
   U6124 : IVI port map( A => n1974, Z => n4950);
   U6125 : IVI port map( A => n288, Z => n4951);
   U6126 : IVI port map( A => n1976, Z => n4952);
   U6127 : IVI port map( A => v_KEY_COLUMN_20_port, Z => n4953);
   U6128 : IVI port map( A => v_KEY_COLUMN_1_port, Z => n4954);
   U6129 : IVI port map( A => n120, Z => n4955);
   U6130 : IVI port map( A => n126, Z => n4956);
   U6131 : IVI port map( A => n189, Z => n4957);
   U6132 : IVI port map( A => v_KEY_COLUMN_15_port, Z => n4958);
   U6133 : IVI port map( A => n403, Z => n4959);
   U6134 : IVI port map( A => n408, Z => n4960);
   U6135 : IVI port map( A => n413, Z => n4961);
   U6136 : IVI port map( A => n420, Z => n4962);
   U6137 : IVI port map( A => v_KEY_COLUMN_12_port, Z => n4963);
   U6138 : IVI port map( A => n344, Z => n4964);
   U6139 : IVI port map( A => n352, Z => n4965);
   U6140 : IVI port map( A => n360, Z => n4966);
   U6141 : IVI port map( A => n370, Z => n4967);
   U6142 : IVI port map( A => v_KEY_COLUMN_0_port, Z => n4968);
   U6143 : IVI port map( A => n659, Z => n4969);
   U6144 : IVI port map( A => n1369, Z => n4970);
   U6145 : IVI port map( A => n1376, Z => n4971);
   U6146 : IVI port map( A => n1387, Z => n4972);
   U6147 : IVI port map( A => n1397, Z => n4973);
   U6148 : IVI port map( A => n1372, Z => n4974);
   U6149 : IVI port map( A => n1379, Z => n4975);
   U6150 : IVI port map( A => n1390, Z => n4976);
   U6151 : IVI port map( A => n1398, Z => n4977);
   U6152 : IVI port map( A => n1373, Z => n4978);
   U6153 : IVI port map( A => n1381, Z => n4979);
   U6154 : IVI port map( A => n1391, Z => n4980);
   U6155 : IVI port map( A => n1399, Z => n4981);
   U6156 : IVI port map( A => n1374, Z => n4982);
   U6157 : IVI port map( A => n1382, Z => n4983);
   U6158 : IVI port map( A => n1392, Z => n4984);
   U6159 : IVI port map( A => n1400, Z => n4985);
   U6160 : IVI port map( A => n1375, Z => n4986);
   U6161 : IVI port map( A => n1383, Z => n4987);
   U6162 : IVI port map( A => n1394, Z => n4988);
   U6163 : IVI port map( A => n1401, Z => n4989);
   U6164 : IVI port map( A => n1380, Z => n4990);
   U6165 : IVI port map( A => n1384, Z => n4991);
   U6166 : IVI port map( A => n1395, Z => n4992);
   U6167 : IVI port map( A => n1402, Z => n4993);
   U6168 : IVI port map( A => n1365, Z => n4994);
   U6169 : IVI port map( A => n1385, Z => n4995);
   U6170 : IVI port map( A => n1393, Z => n4996);
   U6171 : IVI port map( A => n1396, Z => n4997);
   U6172 : IVI port map( A => DATA_I(0), Z => n4998);
   U6173 : IVI port map( A => VALID_DATA_I, Z => n4999);
   U6174 : IVI port map( A => n1360, Z => n5000);
   U6175 : IVI port map( A => n1445, Z => n5001);
   U6176 : IVI port map( A => n1446, Z => n5002);
   U6177 : IVI port map( A => n163, Z => n5003);
   U6178 : IVI port map( A => n164, Z => n5004);
   U6179 : IVI port map( A => n1439, Z => n5005);
   U6180 : IVI port map( A => n1407, Z => n5006);
   U6181 : IVI port map( A => n1410, Z => n5007);
   U6182 : IVI port map( A => n1411, Z => n5008);
   U6183 : IVI port map( A => n1413, Z => n5009);
   U6184 : IVI port map( A => n1433, Z => n5011);
   U6185 : IVI port map( A => n1440, Z => n5012);
   U6186 : IVI port map( A => n1424, Z => n5013);
   U6187 : IVI port map( A => n103, Z => n5014);
   U6188 : IVI port map( A => n1301, Z => n5015);
   U6189 : IVI port map( A => n1343, Z => n5016);
   U6190 : IVI port map( A => n1478, Z => n5017);
   U6191 : IVI port map( A => n3800, Z => n5018);
   U6192 : IVI port map( A => n1479, Z => n5019);
   U6193 : IVI port map( A => n1342, Z => n5021);
   U6194 : IVI port map( A => n1444, Z => n5022);
   U6195 : IVI port map( A => n3672, Z => n5023);
   U6196 : IVI port map( A => n3804, Z => n5024);
   U6197 : IVI port map( A => n3805, Z => n5025);
   U6198 : IVI port map( A => n1457, Z => n5026);
   U6199 : IVI port map( A => n1458, Z => n5027);
   U6200 : IVI port map( A => n2806, Z => n5028);
   U6201 : IVI port map( A => n2598, Z => n5029);
   U6202 : IVI port map( A => n2785, Z => n5030);
   U6203 : IVI port map( A => n2551, Z => n5031);
   U6204 : IVI port map( A => n2669, Z => n5032);
   U6205 : IVI port map( A => n2632, Z => n5033);
   U6206 : IVI port map( A => n2707, Z => n5034);
   U6207 : IVI port map( A => n2845, Z => n5035);
   U6208 : IVI port map( A => n2628, Z => n5036);
   U6209 : IVI port map( A => n2866, Z => n5037);
   U6210 : IVI port map( A => n2686, Z => n5038);
   U6211 : IVI port map( A => n2832, Z => n5039);
   U6212 : IVI port map( A => n2674, Z => n5040);
   U6213 : IVI port map( A => n2534, Z => n5041);
   U6214 : IVI port map( A => n2869, Z => n5042);
   U6215 : IVI port map( A => n2583, Z => n5043);
   U6216 : IVI port map( A => n2731, Z => n5044);
   U6217 : IVI port map( A => n2520, Z => n5045);
   U6218 : IVI port map( A => n2521, Z => n5046);
   U6219 : IVI port map( A => n2516, Z => n5047);
   U6220 : IVI port map( A => n2532, Z => n5048);
   U6221 : IVI port map( A => n2642, Z => n5049);
   U6222 : IVI port map( A => n2670, Z => n5050);
   U6223 : IVI port map( A => n2796, Z => n5051);
   U6224 : IVI port map( A => n2721, Z => n5052);
   U6225 : IVI port map( A => n2793, Z => n5053);
   U6226 : IVI port map( A => n2574, Z => n5054);
   U6227 : IVI port map( A => n2553, Z => n5055);
   U6228 : IVI port map( A => n2617, Z => n5056);
   U6229 : IVI port map( A => n1930, Z => n5057);
   U6230 : IVI port map( A => n2708, Z => n5058);
   U6231 : IVI port map( A => n2499, Z => n5059);
   U6232 : IVI port map( A => n2668, Z => n5060);
   U6233 : IVI port map( A => n2732, Z => n5061);
   U6234 : IVI port map( A => n1964, Z => n5062);
   U6235 : IVI port map( A => n2541, Z => n5063);
   U6236 : IVI port map( A => n2559, Z => n5064);
   U6237 : IVI port map( A => n3039, Z => n5065);
   U6238 : IVI port map( A => n2322, Z => n5066);
   U6239 : IVI port map( A => n1844, Z => n5067);
   U6240 : IVI port map( A => n2395, Z => n5068);
   U6241 : IVI port map( A => n2238, Z => n5069);
   U6242 : IVI port map( A => n1876, Z => n5070);
   U6243 : IVI port map( A => n2268, Z => n5071);
   U6244 : IVI port map( A => n2182, Z => n5072);
   U6245 : IVI port map( A => n3442, Z => n5073);
   U6246 : IVI port map( A => n2657, Z => n5074);
   U6247 : IVI port map( A => n2582, Z => n5075);
   U6248 : IVI port map( A => n2575, Z => n5076);
   U6249 : IVI port map( A => n2542, Z => n5077);
   U6250 : IVI port map( A => n2752, Z => n5078);
   U6251 : IVI port map( A => n2961, Z => n5079);
   U6252 : IVI port map( A => n3049, Z => n5080);
   U6253 : IVI port map( A => n3082, Z => n5081);
   U6254 : IVI port map( A => n2959, Z => n5082);
   U6255 : IVI port map( A => n3078, Z => n5083);
   U6256 : IVI port map( A => n3206, Z => n5084);
   U6257 : IVI port map( A => n3284, Z => n5085);
   U6258 : IVI port map( A => n3281, Z => n5086);
   U6259 : IVI port map( A => n2982, Z => n5087);
   U6260 : IVI port map( A => n2949, Z => n5088);
   U6261 : IVI port map( A => n2966, Z => n5089);
   U6262 : IVI port map( A => n3216, Z => n5090);
   U6263 : IVI port map( A => n3127, Z => n5091);
   U6264 : IVI port map( A => n3195, Z => n5092);
   U6265 : IVI port map( A => n3094, Z => n5093);
   U6266 : IVI port map( A => n3237, Z => n5094);
   U6267 : IVI port map( A => n2989, Z => n5095);
   U6268 : IVI port map( A => n3114, Z => n5096);
   U6269 : IVI port map( A => n3065, Z => n5097);
   U6270 : IVI port map( A => n3203, Z => n5098);
   U6271 : IVI port map( A => n2924, Z => n5099);
   U6272 : IVI port map( A => n1657, Z => n5100);
   U6273 : IVI port map( A => n1694, Z => n5101);
   U6274 : IVI port map( A => n2943, Z => n5102);
   U6275 : IVI port map( A => n1685, Z => n5103);
   U6276 : IVI port map( A => n3137, Z => n5104);
   U6277 : IVI port map( A => n3138, Z => n5105);
   U6278 : IVI port map( A => n3250, Z => n5106);
   U6279 : IVI port map( A => n3005, Z => n5107);
   U6280 : IVI port map( A => n2950, Z => n5108);
   U6281 : IVI port map( A => n3113, Z => n5109);
   U6282 : IVI port map( A => n2981, Z => n5110);
   U6283 : IVI port map( A => n3035, Z => n5111);
   U6284 : IVI port map( A => n3003, Z => n5112);
   U6285 : IVI port map( A => n3159, Z => n5113);
   U6286 : IVI port map( A => n3076, Z => n5114);
   U6287 : IVI port map( A => n2928, Z => n5115);
   U6288 : IVI port map( A => n2231, Z => n5116);
   U6289 : IVI port map( A => n2073, Z => n5117);
   U6290 : IVI port map( A => n1884, Z => n5118);
   U6291 : IVI port map( A => n2148, Z => n5119);
   U6292 : IVI port map( A => n2291, Z => n5120);
   U6293 : IVI port map( A => n2108, Z => n5121);
   U6294 : IVI port map( A => n2144, Z => n5122);
   U6295 : IVI port map( A => n2033, Z => n5123);
   U6296 : IVI port map( A => n2407, Z => n5124);
   U6297 : IVI port map( A => n2394, Z => n5125);
   U6298 : IVI port map( A => n2120, Z => n5126);
   U6299 : IVI port map( A => n2298, Z => n5127);
   U6300 : IVI port map( A => n1892, Z => n5128);
   U6301 : IVI port map( A => n2050, Z => n5129);
   U6302 : IVI port map( A => n2068, Z => n5130);
   U6303 : IVI port map( A => n2316, Z => n5131);
   U6304 : IVI port map( A => n2191, Z => n5132);
   U6305 : IVI port map( A => n2015, Z => n5133);
   U6306 : IVI port map( A => n2093, Z => n5134);
   U6307 : IVI port map( A => n2251, Z => n5135);
   U6308 : IVI port map( A => n1889, Z => n5136);
   U6309 : IVI port map( A => n2168, Z => n5137);
   U6310 : IVI port map( A => n1852, Z => n5138);
   U6311 : IVI port map( A => n2143, Z => n5139);
   U6312 : IVI port map( A => n2021, Z => n5140);
   U6313 : IVI port map( A => n1854, Z => n5141);
   U6314 : IVI port map( A => n1888, Z => n5142);
   U6315 : IVI port map( A => n2216, Z => n5143);
   U6316 : IVI port map( A => n2129, Z => n5144);
   U6317 : IVI port map( A => n2273, Z => n5145);
   U6318 : IVI port map( A => n2071, Z => n5146);
   U6319 : IVI port map( A => n2069, Z => n5147);
   U6320 : IVI port map( A => n2164, Z => n5148);
   U6321 : IVI port map( A => n2095, Z => n5149);
   U6322 : IVI port map( A => n2057, Z => n5150);
   U6323 : IVI port map( A => n2140, Z => n5151);
   U6324 : IVI port map( A => n2032, Z => n5152);
   U6325 : IVI port map( A => n2162, Z => n5153);
   U6326 : IVI port map( A => n2241, Z => n5154);
   U6327 : IVI port map( A => n2214, Z => n5155);
   U6328 : IVI port map( A => n3364, Z => n5156);
   U6329 : IVI port map( A => n3452, Z => n5157);
   U6330 : IVI port map( A => n3485, Z => n5158);
   U6331 : IVI port map( A => n3362, Z => n5159);
   U6332 : IVI port map( A => n3481, Z => n5160);
   U6333 : IVI port map( A => n3610, Z => n5161);
   U6334 : IVI port map( A => n3692, Z => n5162);
   U6335 : IVI port map( A => n3689, Z => n5163);
   U6336 : IVI port map( A => n3385, Z => n5164);
   U6337 : IVI port map( A => n3352, Z => n5165);
   U6338 : IVI port map( A => n3369, Z => n5166);
   U6339 : IVI port map( A => n3620, Z => n5167);
   U6340 : IVI port map( A => n3531, Z => n5168);
   U6341 : IVI port map( A => n3599, Z => n5169);
   U6342 : IVI port map( A => n3497, Z => n5170);
   U6343 : IVI port map( A => n3642, Z => n5171);
   U6344 : IVI port map( A => n3392, Z => n5172);
   U6345 : IVI port map( A => n3518, Z => n5173);
   U6346 : IVI port map( A => n3468, Z => n5174);
   U6347 : IVI port map( A => n3607, Z => n5175);
   U6348 : IVI port map( A => n3327, Z => n5176);
   U6349 : IVI port map( A => n2446, Z => n5177);
   U6350 : IVI port map( A => n2479, Z => n5178);
   U6351 : IVI port map( A => n3346, Z => n5179);
   U6352 : IVI port map( A => n2470, Z => n5180);
   U6353 : IVI port map( A => n3541, Z => n5181);
   U6354 : IVI port map( A => n3542, Z => n5182);
   U6355 : IVI port map( A => n3655, Z => n5183);
   U6356 : IVI port map( A => n3408, Z => n5184);
   U6357 : IVI port map( A => n3353, Z => n5185);
   U6358 : IVI port map( A => n3517, Z => n5186);
   U6359 : IVI port map( A => n3384, Z => n5187);
   U6360 : IVI port map( A => n3438, Z => n5188);
   U6361 : IVI port map( A => n3406, Z => n5189);
   U6362 : IVI port map( A => n3563, Z => n5190);
   U6363 : IVI port map( A => n3479, Z => n5191);
   U6364 : IVI port map( A => n3331, Z => n5192);
   U6365 : IVI port map( A => n2942, Z => n5193);
   U6366 : IVI port map( A => n2945, Z => n5194);
   U6367 : IVI port map( A => n1857, Z => n5195);
   U6368 : IVI port map( A => n2066, Z => n5200);
   U6369 : IVI port map( A => n2116, Z => n5201);
   U6370 : IVI port map( A => n2065, Z => n5202);
   U6371 : IVI port map( A => n2533, Z => n5204);
   U6372 : IVI port map( A => n2536, Z => n5205);
   U6373 : IVI port map( A => n3345, Z => n5206);
   U6374 : IVI port map( A => n3348, Z => n5207);
   U6375 : IVI port map( A => n3387, Z => n5208);
   U6376 : IVI port map( A => n2469, Z => n5209);
   U6377 : IVI port map( A => n3339, Z => n5210);
   U6378 : IVI port map( A => n3321, Z => n5212);
   U6379 : IVI port map( A => n3334, Z => n5213);
   U6380 : IVI port map( A => n3388, Z => n5215);
   U6381 : IVI port map( A => n3454, Z => n5216);
   U6382 : IVI port map( A => n2984, Z => n5217);
   U6383 : IVI port map( A => n1684, Z => n5218);
   U6384 : IVI port map( A => n2936, Z => n5219);
   U6385 : IVI port map( A => n2918, Z => n5221);
   U6386 : IVI port map( A => n2931, Z => n5222);
   U6387 : IVI port map( A => n2985, Z => n5224);
   U6388 : IVI port map( A => n3051, Z => n5225);
   U6389 : IVI port map( A => n2577, Z => n5226);
   U6390 : IVI port map( A => n1954, Z => n5227);
   U6391 : IVI port map( A => n2578, Z => n5228);
   U6392 : IVI port map( A => n2644, Z => n5229);
   U6393 : IVI port map( A => n2526, Z => n5230);
   U6394 : IVI port map( A => n2511, Z => n5232);
   U6395 : IVI port map( A => n2522, Z => n5233);
   U6396 : IVI port map( A => n1881, Z => n5235);
   U6397 : IVI port map( A => n2930, Z => n5236);
   U6398 : IVI port map( A => n2906, Z => n5237);
   U6399 : IVI port map( A => n3077, Z => n5238);
   U6400 : IVI port map( A => n3023, Z => n5239);
   U6401 : IVI port map( A => n2275, Z => n5240);
   U6402 : IVI port map( A => n2072, Z => n5241);
   U6403 : IVI port map( A => n2112, Z => n5242);
   U6404 : IVI port map( A => n3333, Z => n5243);
   U6405 : IVI port map( A => n3309, Z => n5244);
   U6406 : IVI port map( A => n3480, Z => n5245);
   U6407 : IVI port map( A => n3426, Z => n5246);

end SYN_Behavioral;
