
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_aes_dec_KEY_SIZE2 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_aes_dec_KEY_SIZE2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_aes_dec_KEY_SIZE2.all;

entity key_expansion is

   port( KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, CLK_I, RESET_I
         , CE_I : in std_logic;  DONE_O : out std_logic;  GET_KEY_I : in 
         std_logic;  KEY_NUMB_I : in std_logic_vector (5 downto 0);  KEY_EXP_O 
         : out std_logic_vector (31 downto 0));

end key_expansion;

architecture SYN_Behavioral of key_expansion is

   component NR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component IV
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21L
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AN2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component NR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AN3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EON1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO7
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX31L
      port( D0, D1, D2, A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EO
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21H
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EN
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FD1
      port( D, CP : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal v_KEY32_IN_31_port, v_KEY32_IN_30_port, v_KEY32_IN_29_port, 
      v_KEY32_IN_28_port, v_KEY32_IN_27_port, v_KEY32_IN_26_port, 
      v_KEY32_IN_25_port, v_KEY32_IN_24_port, v_KEY32_IN_23_port, 
      v_KEY32_IN_22_port, v_KEY32_IN_21_port, v_KEY32_IN_20_port, 
      v_KEY32_IN_19_port, v_KEY32_IN_18_port, v_KEY32_IN_17_port, 
      v_KEY32_IN_16_port, v_KEY32_IN_15_port, v_KEY32_IN_14_port, 
      v_KEY32_IN_13_port, v_KEY32_IN_12_port, v_KEY32_IN_11_port, 
      v_KEY32_IN_10_port, v_KEY32_IN_9_port, v_KEY32_IN_8_port, 
      v_KEY32_IN_7_port, v_KEY32_IN_6_port, v_KEY32_IN_5_port, 
      v_KEY32_IN_4_port, v_KEY32_IN_3_port, v_KEY32_IN_2_port, 
      v_KEY32_IN_1_port, v_KEY32_IN_0_port, v_CALCULATION_CNTR_7_port, 
      v_CALCULATION_CNTR_6_port, v_CALCULATION_CNTR_5_port, 
      v_CALCULATION_CNTR_4_port, v_CALCULATION_CNTR_3_port, 
      v_CALCULATION_CNTR_2_port, v_CALCULATION_CNTR_1_port, 
      v_CALCULATION_CNTR_0_port, v_KEY_COL_OUT0_31_port, v_KEY_COL_OUT0_30_port
      , v_KEY_COL_OUT0_29_port, v_KEY_COL_OUT0_28_port, v_KEY_COL_OUT0_27_port,
      v_KEY_COL_OUT0_26_port, v_KEY_COL_OUT0_25_port, v_KEY_COL_OUT0_24_port, 
      v_KEY_COL_OUT0_23_port, v_KEY_COL_OUT0_22_port, v_KEY_COL_OUT0_21_port, 
      v_KEY_COL_OUT0_20_port, v_KEY_COL_OUT0_19_port, v_KEY_COL_OUT0_18_port, 
      v_KEY_COL_OUT0_17_port, v_KEY_COL_OUT0_16_port, v_KEY_COL_OUT0_15_port, 
      v_KEY_COL_OUT0_14_port, v_KEY_COL_OUT0_13_port, v_KEY_COL_OUT0_12_port, 
      v_KEY_COL_OUT0_11_port, v_KEY_COL_OUT0_10_port, v_KEY_COL_OUT0_9_port, 
      v_KEY_COL_OUT0_8_port, v_KEY_COL_OUT0_5_port, v_KEY_COL_OUT0_4_port, 
      v_KEY_COL_OUT0_3_port, v_KEY_COL_OUT0_2_port, v_KEY_COL_OUT0_1_port, 
      v_TEMP_VECTOR_31_port, v_TEMP_VECTOR_30_port, v_TEMP_VECTOR_29_port, 
      v_TEMP_VECTOR_28_port, v_TEMP_VECTOR_27_port, v_TEMP_VECTOR_26_port, 
      v_TEMP_VECTOR_25_port, v_TEMP_VECTOR_24_port, v_TEMP_VECTOR_23_port, 
      v_TEMP_VECTOR_22_port, v_TEMP_VECTOR_21_port, v_TEMP_VECTOR_20_port, 
      v_TEMP_VECTOR_19_port, v_TEMP_VECTOR_18_port, v_TEMP_VECTOR_17_port, 
      v_TEMP_VECTOR_16_port, v_TEMP_VECTOR_15_port, v_TEMP_VECTOR_14_port, 
      v_TEMP_VECTOR_13_port, v_TEMP_VECTOR_12_port, v_TEMP_VECTOR_11_port, 
      v_TEMP_VECTOR_10_port, v_TEMP_VECTOR_9_port, v_TEMP_VECTOR_8_port, 
      v_TEMP_VECTOR_7_port, v_TEMP_VECTOR_6_port, v_TEMP_VECTOR_5_port, 
      v_TEMP_VECTOR_4_port, v_TEMP_VECTOR_3_port, v_TEMP_VECTOR_2_port, 
      v_TEMP_VECTOR_1_port, v_TEMP_VECTOR_0_port, v_SUB_WORD_7_port, 
      v_SUB_WORD_6_port, v_SUB_WORD_0_port, n2489, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
      n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, 
      n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
      n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
      n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
      n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
      n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, 
      n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, 
      n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
      n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, 
      n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, 
      n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
      n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, 
      n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, 
      n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
      n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
      n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
      n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
      n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
      n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, 
      n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, 
      n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, 
      n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, 
      n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, 
      n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, 
      n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, 
      n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, 
      n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, 
      n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, 
      n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, 
      n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, 
      n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, 
      n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, 
      n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, 
      n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, 
      n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
      n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, 
      n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, 
      n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, 
      n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, 
      n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, 
      n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, 
      n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, 
      n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, 
      n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, 
      n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, 
      n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, 
      n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, 
      n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, 
      n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, 
      n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, 
      n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, 
      n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, 
      n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, 
      n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, 
      n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, 
      n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, 
      n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, 
      n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, 
      n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, 
      n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, 
      n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, 
      n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, 
      n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, 
      n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, 
      n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, 
      n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, 
      n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, 
      n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, 
      n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, 
      n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, 
      n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, 
      n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, 
      n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, 
      n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
      n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, 
      n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, 
      n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, 
      n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
      n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, 
      n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, 
      n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
      n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, 
      n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, 
      n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, 
      n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, 
      n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, 
      n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, 
      n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, 
      n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, 
      n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, 
      n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, 
      n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, 
      n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, 
      n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, 
      n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, 
      n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, 
      n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, 
      n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, 
      n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, 
      n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, 
      n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, 
      n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, 
      n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, 
      n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, 
      n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, 
      n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, 
      n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, 
      n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, 
      n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, 
      n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, 
      n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, 
      n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, 
      n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, 
      n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, 
      n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, 
      n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, 
      n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, 
      n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, 
      n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, 
      n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, 
      n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, 
      n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, 
      n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, 
      n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, 
      n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, 
      n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, 
      n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, 
      n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, 
      n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, 
      n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, 
      n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, 
      n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, 
      n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, 
      n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, 
      n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, 
      n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, 
      n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, 
      n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, 
      n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, 
      n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, 
      n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, 
      n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, 
      n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, 
      n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, 
      n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, 
      n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, 
      n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, 
      n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, 
      n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, 
      n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, 
      n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, 
      n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, 
      n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, 
      n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, 
      n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, 
      n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, 
      n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, 
      n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, 
      n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6651, n6652, n6653, 
      n6654, n6655, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, 
      n6712, n6713, n6714, n6715, n6748, n6749, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, 
      n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, 
      n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, 
      n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, 
      n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
      n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, 
      n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, 
      n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
      n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, 
      n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
      n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, 
      n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, 
      n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
      n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
      n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
      n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, 
      n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
      n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, 
      n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, 
      n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, 
      n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
      n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, 
      n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
      n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
      n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
      n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, 
      n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
      n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
      n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, 
      n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
      n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, 
      n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, 
      n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, 
      n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
      n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
      n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, 
      n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, 
      n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, 
      n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
      n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, 
      n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, 
      n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, 
      n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, 
      n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, 
      n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, 
      n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, 
      n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, 
      n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, 
      n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, 
      n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, 
      n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, 
      n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
      n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
      n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
      n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, 
      n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
      n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
      n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
      n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, 
      n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, 
      n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, 
      n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, 
      n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
      n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, 
      n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, 
      n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, 
      n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, 
      n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, 
      n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, 
      n2488, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
      n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, 
      n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, 
      n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, 
      n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, 
      n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
      n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, 
      n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, 
      n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, 
      n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
      n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
      n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, 
      n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, 
      n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
      n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, 
      n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, 
      n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
      n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
      n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
      n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
      n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
      n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
      n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
      n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, 
      n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
      n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
      n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
      n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
      n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
      n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
      n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
      n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
      n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, 
      n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
      n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
      n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
      n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, 
      n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
      n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, 
      n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
      n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
      n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, 
      n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
      n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, 
      n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
      n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, 
      n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
      n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, 
      n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
      n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, 
      n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, 
      n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, 
      n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, 
      n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, 
      n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, 
      n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, 
      n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, 
      n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, 
      n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, 
      n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, 
      n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, 
      n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, 
      n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, 
      n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, 
      n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, 
      n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, 
      n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, 
      n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, 
      n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, 
      n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, 
      n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, 
      n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, 
      n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
      n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, 
      n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
      n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, 
      n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, 
      n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, 
      n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
      n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, 
      n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, 
      n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, 
      n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
      n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, 
      n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
      n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, 
      n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
      n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, 
      n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
      n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
      n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
      n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, 
      n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
      n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, 
      n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
      n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, 
      n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
      n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, 
      n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, 
      n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, 
      n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, 
      n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, 
      n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, 
      n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, 
      n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, 
      n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, 
      n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, 
      n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, 
      n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, 
      n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, 
      n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, 
      n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, 
      n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
      n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, 
      n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, 
      n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
      n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, 
      n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, 
      n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, 
      n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, 
      n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
      n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, 
      n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, 
      n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
      n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
      n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n_1000, n_1001, 
      n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, 
      n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, 
      n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, 
      n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, 
      n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, 
      n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, 
      n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, 
      n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, 
      n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, 
      n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, 
      n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, 
      n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, 
      n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, 
      n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, 
      n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, 
      n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, 
      n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, 
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, 
      n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, 
      n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, 
      n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, 
      n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, 
      n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, 
      n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, 
      n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, 
      n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, 
      n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, 
      n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, 
      n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, 
      n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, 
      n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, 
      n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, 
      n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, 
      n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, 
      n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, 
      n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, 
      n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, 
      n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, 
      n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, 
      n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, 
      n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, 
      n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, 
      n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, 
      n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, 
      n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, 
      n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, 
      n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, 
      n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, 
      n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, 
      n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, 
      n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, 
      n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, 
      n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, 
      n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, 
      n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, 
      n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, 
      n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, 
      n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, 
      n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, 
      n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, 
      n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, 
      n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, 
      n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, 
      n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, 
      n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, 
      n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, 
      n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, 
      n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, 
      n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, 
      n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, 
      n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, 
      n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, 
      n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, 
      n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, 
      n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, 
      n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, 
      n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, 
      n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, 
      n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, 
      n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, 
      n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, 
      n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, 
      n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, 
      n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, 
      n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, 
      n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, 
      n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, 
      n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, 
      n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, 
      n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, 
      n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, 
      n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, 
      n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, 
      n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, 
      n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, 
      n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, 
      n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, 
      n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, 
      n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, 
      n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, 
      n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, 
      n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, 
      n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, 
      n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, 
      n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, 
      n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, 
      n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, 
      n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, 
      n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, 
      n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, 
      n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, 
      n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, 
      n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, 
      n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, 
      n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, 
      n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, 
      n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, 
      n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, 
      n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, 
      n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, 
      n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, 
      n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, 
      n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, 
      n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, 
      n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, 
      n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, 
      n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, 
      n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, 
      n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, 
      n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, 
      n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, 
      n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, 
      n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, 
      n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, 
      n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, 
      n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, 
      n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, 
      n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, 
      n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, 
      n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, 
      n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, 
      n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, 
      n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, 
      n_3108, n_3109, n_3110, n_3111 : std_logic;

begin
   
   i_BYTE_CNTR4_reg_0_inst : FD1 port map( D => n6749, CP => CLK_I, Q => n4464,
                           QN => n1039);
   i_BYTE_CNTR4_reg_1_inst : FD1 port map( D => n6748, CP => CLK_I, Q => n4463,
                           QN => n6);
   FF_VALID_KEY_reg : FD1 port map( D => n4589, CP => CLK_I, Q => n4469, QN => 
                           n1040);
   v_KEY32_IN_reg_31_inst : FD1 port map( D => n4479, CP => CLK_I, Q => 
                           v_KEY32_IN_31_port, QN => n_1000);
   v_KEY32_IN_reg_30_inst : FD1 port map( D => n4478, CP => CLK_I, Q => 
                           v_KEY32_IN_30_port, QN => n_1001);
   v_KEY32_IN_reg_29_inst : FD1 port map( D => n4477, CP => CLK_I, Q => 
                           v_KEY32_IN_29_port, QN => n_1002);
   v_KEY32_IN_reg_28_inst : FD1 port map( D => n4476, CP => CLK_I, Q => 
                           v_KEY32_IN_28_port, QN => n_1003);
   v_KEY32_IN_reg_27_inst : FD1 port map( D => n4475, CP => CLK_I, Q => 
                           v_KEY32_IN_27_port, QN => n_1004);
   v_KEY32_IN_reg_26_inst : FD1 port map( D => n4474, CP => CLK_I, Q => 
                           v_KEY32_IN_26_port, QN => n_1005);
   v_KEY32_IN_reg_25_inst : FD1 port map( D => n4473, CP => CLK_I, Q => 
                           v_KEY32_IN_25_port, QN => n_1006);
   v_KEY32_IN_reg_24_inst : FD1 port map( D => n4472, CP => CLK_I, Q => 
                           v_KEY32_IN_24_port, QN => n_1007);
   v_KEY32_IN_reg_23_inst : FD1 port map( D => n4495, CP => CLK_I, Q => 
                           v_KEY32_IN_23_port, QN => n_1008);
   v_KEY32_IN_reg_22_inst : FD1 port map( D => n4494, CP => CLK_I, Q => 
                           v_KEY32_IN_22_port, QN => n_1009);
   v_KEY32_IN_reg_21_inst : FD1 port map( D => n4493, CP => CLK_I, Q => 
                           v_KEY32_IN_21_port, QN => n_1010);
   v_KEY32_IN_reg_20_inst : FD1 port map( D => n4492, CP => CLK_I, Q => 
                           v_KEY32_IN_20_port, QN => n_1011);
   v_KEY32_IN_reg_19_inst : FD1 port map( D => n4491, CP => CLK_I, Q => 
                           v_KEY32_IN_19_port, QN => n_1012);
   v_KEY32_IN_reg_18_inst : FD1 port map( D => n4490, CP => CLK_I, Q => 
                           v_KEY32_IN_18_port, QN => n_1013);
   v_KEY32_IN_reg_17_inst : FD1 port map( D => n4489, CP => CLK_I, Q => 
                           v_KEY32_IN_17_port, QN => n_1014);
   v_KEY32_IN_reg_16_inst : FD1 port map( D => n4488, CP => CLK_I, Q => 
                           v_KEY32_IN_16_port, QN => n_1015);
   v_KEY32_IN_reg_15_inst : FD1 port map( D => n4503, CP => CLK_I, Q => 
                           v_KEY32_IN_15_port, QN => n_1016);
   v_KEY32_IN_reg_14_inst : FD1 port map( D => n4502, CP => CLK_I, Q => 
                           v_KEY32_IN_14_port, QN => n_1017);
   v_KEY32_IN_reg_13_inst : FD1 port map( D => n4501, CP => CLK_I, Q => 
                           v_KEY32_IN_13_port, QN => n_1018);
   v_KEY32_IN_reg_12_inst : FD1 port map( D => n4500, CP => CLK_I, Q => 
                           v_KEY32_IN_12_port, QN => n_1019);
   v_KEY32_IN_reg_11_inst : FD1 port map( D => n4499, CP => CLK_I, Q => 
                           v_KEY32_IN_11_port, QN => n_1020);
   v_KEY32_IN_reg_10_inst : FD1 port map( D => n4498, CP => CLK_I, Q => 
                           v_KEY32_IN_10_port, QN => n_1021);
   v_KEY32_IN_reg_9_inst : FD1 port map( D => n4497, CP => CLK_I, Q => 
                           v_KEY32_IN_9_port, QN => n_1022);
   v_KEY32_IN_reg_8_inst : FD1 port map( D => n4496, CP => CLK_I, Q => 
                           v_KEY32_IN_8_port, QN => n_1023);
   v_KEY32_IN_reg_7_inst : FD1 port map( D => n4487, CP => CLK_I, Q => 
                           v_KEY32_IN_7_port, QN => n2119);
   v_KEY32_IN_reg_6_inst : FD1 port map( D => n4486, CP => CLK_I, Q => 
                           v_KEY32_IN_6_port, QN => n2117);
   v_KEY32_IN_reg_5_inst : FD1 port map( D => n4485, CP => CLK_I, Q => 
                           v_KEY32_IN_5_port, QN => n2116);
   v_KEY32_IN_reg_4_inst : FD1 port map( D => n4484, CP => CLK_I, Q => 
                           v_KEY32_IN_4_port, QN => n2115);
   v_KEY32_IN_reg_3_inst : FD1 port map( D => n4483, CP => CLK_I, Q => 
                           v_KEY32_IN_3_port, QN => n2114);
   v_KEY32_IN_reg_2_inst : FD1 port map( D => n4482, CP => CLK_I, Q => 
                           v_KEY32_IN_2_port, QN => n2112);
   v_KEY32_IN_reg_1_inst : FD1 port map( D => n4481, CP => CLK_I, Q => 
                           v_KEY32_IN_1_port, QN => n2111);
   v_KEY32_IN_reg_0_inst : FD1 port map( D => n4480, CP => CLK_I, Q => 
                           v_KEY32_IN_0_port, QN => n2109);
   FF_GET_KEY_reg : FD1 port map( D => GET_KEY_I, CP => CLK_I, Q => n_1024, QN 
                           => n1034);
   v_SUB_WORD_reg_7_inst : FD1 port map( D => n4588, CP => CLK_I, Q => 
                           v_SUB_WORD_7_port, QN => n1075);
   v_SUB_WORD_reg_6_inst : FD1 port map( D => n4587, CP => CLK_I, Q => 
                           v_SUB_WORD_6_port, QN => n1041);
   v_SUB_WORD_reg_5_inst : FD1 port map( D => n4586, CP => CLK_I, Q => n2105, 
                           QN => n4468);
   v_SUB_WORD_reg_4_inst : FD1 port map( D => n4585, CP => CLK_I, Q => n2106, 
                           QN => n4467);
   v_SUB_WORD_reg_3_inst : FD1 port map( D => n4584, CP => CLK_I, Q => n2107, 
                           QN => n4466);
   v_SUB_WORD_reg_2_inst : FD1 port map( D => n4583, CP => CLK_I, Q => n2113, 
                           QN => n4465);
   v_SUB_WORD_reg_1_inst : FD1 port map( D => n4582, CP => CLK_I, Q => n2108, 
                           QN => n4456);
   v_SUB_WORD_reg_0_inst : FD1 port map( D => n4581, CP => CLK_I, Q => 
                           v_SUB_WORD_0_port, QN => n1074);
   v_CALCULATION_CNTR_reg_0_inst : FD1 port map( D => n6651, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_0_port, QN => n1077);
   i_ROUND_reg_3_inst : FD1 port map( D => n6715, CP => CLK_I, Q => n4462, QN 
                           => n1042);
   START_CALCULATION_reg : FD1 port map( D => n6711, CP => CLK_I, Q => n4471, 
                           QN => n1043);
   i_ROUND_reg_0_inst : FD1 port map( D => n6714, CP => CLK_I, Q => n4461, QN 
                           => n3);
   i_ROUND_reg_1_inst : FD1 port map( D => n6713, CP => CLK_I, Q => n4460, QN 
                           => n2104);
   i_ROUND_reg_2_inst : FD1 port map( D => n6712, CP => CLK_I, Q => n4458, QN 
                           => n5);
   DONE_O_reg : FD1 port map( D => n6710, CP => CLK_I, Q => DONE_O, QN => n2489
                           );
   CALCULATION_reg : FD1 port map( D => n6709, CP => CLK_I, Q => n_1025, QN => 
                           n4455);
   v_CALCULATION_CNTR_reg_1_inst : FD1 port map( D => n6652, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_1_port, QN => n7);
   v_CALCULATION_CNTR_reg_2_inst : FD1 port map( D => n6653, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_2_port, QN => n1036);
   v_CALCULATION_CNTR_reg_3_inst : FD1 port map( D => n6654, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_3_port, QN => n1078);
   v_CALCULATION_CNTR_reg_4_inst : FD1 port map( D => n6655, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_4_port, QN => n8);
   v_CALCULATION_CNTR_reg_5_inst : FD1 port map( D => n4504, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_5_port, QN => n_1026);
   v_CALCULATION_CNTR_reg_6_inst : FD1 port map( D => n4505, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_6_port, QN => n1079);
   v_CALCULATION_CNTR_reg_7_inst : FD1 port map( D => n4506, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_7_port, QN => n_1027);
   i_INTERN_ADDR_RD0_reg_0_inst : FD1 port map( D => n6708, CP => CLK_I, Q => 
                           n1, QN => n6649);
   i_INTERN_ADDR_RD0_reg_1_inst : FD1 port map( D => n6707, CP => CLK_I, Q => 
                           n1033, QN => n6648);
   i_INTERN_ADDR_RD0_reg_2_inst : FD1 port map( D => n6706, CP => CLK_I, Q => 
                           n_1028, QN => n6647);
   i_INTERN_ADDR_RD0_reg_3_inst : FD1 port map( D => n6705, CP => CLK_I, Q => 
                           n1044, QN => n6646);
   i_INTERN_ADDR_RD0_reg_4_inst : FD1 port map( D => n6704, CP => CLK_I, Q => 
                           n1037, QN => n6645);
   i_INTERN_ADDR_RD0_reg_5_inst : FD1 port map( D => n6703, CP => CLK_I, Q => 
                           n_1029, QN => n6644);
   SRAM_WREN0_reg : FD1 port map( D => n6702, CP => CLK_I, Q => n4470, QN => 
                           n1076);
   i_SRAM_ADDR_WR0_reg_5_inst : FD1 port map( D => n6701, CP => CLK_I, Q => 
                           n_1030, QN => n6638);
   i_SRAM_ADDR_WR0_reg_0_inst : FD1 port map( D => n6700, CP => CLK_I, Q => n4,
                           QN => n6643);
   i_SRAM_ADDR_WR0_reg_1_inst : FD1 port map( D => n6699, CP => CLK_I, Q => 
                           n1038, QN => n6642);
   i_SRAM_ADDR_WR0_reg_2_inst : FD1 port map( D => n6698, CP => CLK_I, Q => 
                           n_1031, QN => n6641);
   i_SRAM_ADDR_WR0_reg_3_inst : FD1 port map( D => n6697, CP => CLK_I, Q => 
                           n1035, QN => n6640);
   i_SRAM_ADDR_WR0_reg_4_inst : FD1 port map( D => n6696, CP => CLK_I, Q => n2,
                           QN => n6639);
   v_TEMP_VECTOR_reg_7_inst : FD1 port map( D => n6688, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_7_port, QN => n_1032);
   KEY_EXPAN0_reg_63_7_inst : FD1 port map( D => n5101, CP => CLK_I, Q => 
                           n_1033, QN => n1099);
   KEY_EXPAN0_reg_62_7_inst : FD1 port map( D => n5100, CP => CLK_I, Q => 
                           n_1034, QN => n28);
   KEY_EXPAN0_reg_61_7_inst : FD1 port map( D => n5099, CP => CLK_I, Q => 
                           n_1035, QN => n1098);
   KEY_EXPAN0_reg_60_7_inst : FD1 port map( D => n5098, CP => CLK_I, Q => 
                           n_1036, QN => n27);
   KEY_EXPAN0_reg_59_7_inst : FD1 port map( D => n5097, CP => CLK_I, Q => 
                           n_1037, QN => n1097);
   KEY_EXPAN0_reg_58_7_inst : FD1 port map( D => n5096, CP => CLK_I, Q => 
                           n_1038, QN => n26);
   KEY_EXPAN0_reg_57_7_inst : FD1 port map( D => n5095, CP => CLK_I, Q => 
                           n_1039, QN => n1096);
   KEY_EXPAN0_reg_56_7_inst : FD1 port map( D => n5094, CP => CLK_I, Q => 
                           n_1040, QN => n25);
   KEY_EXPAN0_reg_55_7_inst : FD1 port map( D => n5093, CP => CLK_I, Q => 
                           n_1041, QN => n1103);
   KEY_EXPAN0_reg_54_7_inst : FD1 port map( D => n5092, CP => CLK_I, Q => 
                           n_1042, QN => n32);
   KEY_EXPAN0_reg_53_7_inst : FD1 port map( D => n5091, CP => CLK_I, Q => 
                           n_1043, QN => n1102);
   KEY_EXPAN0_reg_52_7_inst : FD1 port map( D => n5090, CP => CLK_I, Q => 
                           n_1044, QN => n31);
   KEY_EXPAN0_reg_51_7_inst : FD1 port map( D => n5089, CP => CLK_I, Q => 
                           n_1045, QN => n1101);
   KEY_EXPAN0_reg_50_7_inst : FD1 port map( D => n5088, CP => CLK_I, Q => 
                           n_1046, QN => n30);
   KEY_EXPAN0_reg_49_7_inst : FD1 port map( D => n5087, CP => CLK_I, Q => 
                           n_1047, QN => n1100);
   KEY_EXPAN0_reg_48_7_inst : FD1 port map( D => n5086, CP => CLK_I, Q => 
                           n_1048, QN => n29);
   KEY_EXPAN0_reg_47_7_inst : FD1 port map( D => n5085, CP => CLK_I, Q => 
                           n_1049, QN => n1107);
   KEY_EXPAN0_reg_46_7_inst : FD1 port map( D => n5084, CP => CLK_I, Q => 
                           n_1050, QN => n36);
   KEY_EXPAN0_reg_45_7_inst : FD1 port map( D => n5083, CP => CLK_I, Q => 
                           n_1051, QN => n1106);
   KEY_EXPAN0_reg_44_7_inst : FD1 port map( D => n5082, CP => CLK_I, Q => 
                           n_1052, QN => n35);
   KEY_EXPAN0_reg_43_7_inst : FD1 port map( D => n5081, CP => CLK_I, Q => 
                           n_1053, QN => n1105);
   KEY_EXPAN0_reg_42_7_inst : FD1 port map( D => n5080, CP => CLK_I, Q => 
                           n_1054, QN => n34);
   KEY_EXPAN0_reg_41_7_inst : FD1 port map( D => n5079, CP => CLK_I, Q => 
                           n_1055, QN => n1104);
   KEY_EXPAN0_reg_40_7_inst : FD1 port map( D => n5078, CP => CLK_I, Q => 
                           n_1056, QN => n33);
   KEY_EXPAN0_reg_39_7_inst : FD1 port map( D => n5077, CP => CLK_I, Q => 
                           n_1057, QN => n1111);
   KEY_EXPAN0_reg_38_7_inst : FD1 port map( D => n5076, CP => CLK_I, Q => 
                           n_1058, QN => n40);
   KEY_EXPAN0_reg_37_7_inst : FD1 port map( D => n5075, CP => CLK_I, Q => 
                           n_1059, QN => n1110);
   KEY_EXPAN0_reg_36_7_inst : FD1 port map( D => n5074, CP => CLK_I, Q => 
                           n_1060, QN => n39);
   KEY_EXPAN0_reg_35_7_inst : FD1 port map( D => n5073, CP => CLK_I, Q => 
                           n_1061, QN => n1109);
   KEY_EXPAN0_reg_34_7_inst : FD1 port map( D => n5072, CP => CLK_I, Q => 
                           n_1062, QN => n38);
   KEY_EXPAN0_reg_33_7_inst : FD1 port map( D => n5071, CP => CLK_I, Q => 
                           n_1063, QN => n1108);
   KEY_EXPAN0_reg_32_7_inst : FD1 port map( D => n5070, CP => CLK_I, Q => 
                           n_1064, QN => n37);
   KEY_EXPAN0_reg_31_7_inst : FD1 port map( D => n5069, CP => CLK_I, Q => 
                           n_1065, QN => n1083);
   KEY_EXPAN0_reg_30_7_inst : FD1 port map( D => n5068, CP => CLK_I, Q => 
                           n_1066, QN => n12);
   KEY_EXPAN0_reg_29_7_inst : FD1 port map( D => n5067, CP => CLK_I, Q => 
                           n_1067, QN => n1082);
   KEY_EXPAN0_reg_28_7_inst : FD1 port map( D => n5066, CP => CLK_I, Q => 
                           n_1068, QN => n11);
   KEY_EXPAN0_reg_27_7_inst : FD1 port map( D => n5065, CP => CLK_I, Q => 
                           n_1069, QN => n1081);
   KEY_EXPAN0_reg_26_7_inst : FD1 port map( D => n5064, CP => CLK_I, Q => 
                           n_1070, QN => n10);
   KEY_EXPAN0_reg_25_7_inst : FD1 port map( D => n5063, CP => CLK_I, Q => 
                           n_1071, QN => n1080);
   KEY_EXPAN0_reg_24_7_inst : FD1 port map( D => n5062, CP => CLK_I, Q => 
                           n_1072, QN => n9);
   KEY_EXPAN0_reg_23_7_inst : FD1 port map( D => n5061, CP => CLK_I, Q => 
                           n_1073, QN => n1087);
   KEY_EXPAN0_reg_22_7_inst : FD1 port map( D => n5060, CP => CLK_I, Q => 
                           n_1074, QN => n16);
   KEY_EXPAN0_reg_21_7_inst : FD1 port map( D => n5059, CP => CLK_I, Q => 
                           n_1075, QN => n1086);
   KEY_EXPAN0_reg_20_7_inst : FD1 port map( D => n5058, CP => CLK_I, Q => 
                           n_1076, QN => n15);
   KEY_EXPAN0_reg_19_7_inst : FD1 port map( D => n5057, CP => CLK_I, Q => 
                           n_1077, QN => n1085);
   KEY_EXPAN0_reg_18_7_inst : FD1 port map( D => n5056, CP => CLK_I, Q => 
                           n_1078, QN => n14);
   KEY_EXPAN0_reg_17_7_inst : FD1 port map( D => n5055, CP => CLK_I, Q => 
                           n_1079, QN => n1084);
   KEY_EXPAN0_reg_16_7_inst : FD1 port map( D => n5054, CP => CLK_I, Q => 
                           n_1080, QN => n13);
   KEY_EXPAN0_reg_15_7_inst : FD1 port map( D => n5053, CP => CLK_I, Q => 
                           n_1081, QN => n1091);
   KEY_EXPAN0_reg_14_7_inst : FD1 port map( D => n5052, CP => CLK_I, Q => 
                           n_1082, QN => n20);
   KEY_EXPAN0_reg_13_7_inst : FD1 port map( D => n5051, CP => CLK_I, Q => 
                           n_1083, QN => n1090);
   KEY_EXPAN0_reg_12_7_inst : FD1 port map( D => n5050, CP => CLK_I, Q => 
                           n_1084, QN => n19);
   KEY_EXPAN0_reg_11_7_inst : FD1 port map( D => n5049, CP => CLK_I, Q => 
                           n_1085, QN => n1089);
   KEY_EXPAN0_reg_10_7_inst : FD1 port map( D => n5048, CP => CLK_I, Q => 
                           n_1086, QN => n18);
   KEY_EXPAN0_reg_9_7_inst : FD1 port map( D => n5047, CP => CLK_I, Q => n_1087
                           , QN => n1088);
   KEY_EXPAN0_reg_8_7_inst : FD1 port map( D => n5046, CP => CLK_I, Q => n_1088
                           , QN => n17);
   KEY_EXPAN0_reg_7_7_inst : FD1 port map( D => n5045, CP => CLK_I, Q => n_1089
                           , QN => n1095);
   KEY_EXPAN0_reg_6_7_inst : FD1 port map( D => n5044, CP => CLK_I, Q => n_1090
                           , QN => n24);
   KEY_EXPAN0_reg_5_7_inst : FD1 port map( D => n5043, CP => CLK_I, Q => n_1091
                           , QN => n1094);
   KEY_EXPAN0_reg_4_7_inst : FD1 port map( D => n5042, CP => CLK_I, Q => n_1092
                           , QN => n23);
   KEY_EXPAN0_reg_3_7_inst : FD1 port map( D => n5041, CP => CLK_I, Q => n_1093
                           , QN => n1093);
   KEY_EXPAN0_reg_2_7_inst : FD1 port map( D => n5040, CP => CLK_I, Q => n_1094
                           , QN => n22);
   KEY_EXPAN0_reg_1_7_inst : FD1 port map( D => n5039, CP => CLK_I, Q => n_1095
                           , QN => n1092);
   KEY_EXPAN0_reg_0_7_inst : FD1 port map( D => n5038, CP => CLK_I, Q => n_1096
                           , QN => n21);
   v_KEY_COL_OUT0_reg_7_inst : FD1 port map( D => n4580, CP => CLK_I, Q => 
                           n2120, QN => n4454);
   v_TEMP_VECTOR_reg_31_inst : FD1 port map( D => n6664, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_31_port, QN => n_1097);
   KEY_EXPAN0_reg_63_31_inst : FD1 port map( D => n6637, CP => CLK_I, Q => 
                           n_1098, QN => n1131);
   KEY_EXPAN0_reg_62_31_inst : FD1 port map( D => n6636, CP => CLK_I, Q => 
                           n_1099, QN => n60);
   KEY_EXPAN0_reg_61_31_inst : FD1 port map( D => n6635, CP => CLK_I, Q => 
                           n_1100, QN => n1130);
   KEY_EXPAN0_reg_60_31_inst : FD1 port map( D => n6634, CP => CLK_I, Q => 
                           n_1101, QN => n59);
   KEY_EXPAN0_reg_59_31_inst : FD1 port map( D => n6633, CP => CLK_I, Q => 
                           n_1102, QN => n1129);
   KEY_EXPAN0_reg_58_31_inst : FD1 port map( D => n6632, CP => CLK_I, Q => 
                           n_1103, QN => n58);
   KEY_EXPAN0_reg_57_31_inst : FD1 port map( D => n6631, CP => CLK_I, Q => 
                           n_1104, QN => n1128);
   KEY_EXPAN0_reg_56_31_inst : FD1 port map( D => n6630, CP => CLK_I, Q => 
                           n_1105, QN => n57);
   KEY_EXPAN0_reg_55_31_inst : FD1 port map( D => n6629, CP => CLK_I, Q => 
                           n_1106, QN => n1135);
   KEY_EXPAN0_reg_54_31_inst : FD1 port map( D => n6628, CP => CLK_I, Q => 
                           n_1107, QN => n64);
   KEY_EXPAN0_reg_53_31_inst : FD1 port map( D => n6627, CP => CLK_I, Q => 
                           n_1108, QN => n1134);
   KEY_EXPAN0_reg_52_31_inst : FD1 port map( D => n6626, CP => CLK_I, Q => 
                           n_1109, QN => n63);
   KEY_EXPAN0_reg_51_31_inst : FD1 port map( D => n6625, CP => CLK_I, Q => 
                           n_1110, QN => n1133);
   KEY_EXPAN0_reg_50_31_inst : FD1 port map( D => n6624, CP => CLK_I, Q => 
                           n_1111, QN => n62);
   KEY_EXPAN0_reg_49_31_inst : FD1 port map( D => n6623, CP => CLK_I, Q => 
                           n_1112, QN => n1132);
   KEY_EXPAN0_reg_48_31_inst : FD1 port map( D => n6622, CP => CLK_I, Q => 
                           n_1113, QN => n61);
   KEY_EXPAN0_reg_47_31_inst : FD1 port map( D => n6621, CP => CLK_I, Q => 
                           n_1114, QN => n1139);
   KEY_EXPAN0_reg_46_31_inst : FD1 port map( D => n6620, CP => CLK_I, Q => 
                           n_1115, QN => n68);
   KEY_EXPAN0_reg_45_31_inst : FD1 port map( D => n6619, CP => CLK_I, Q => 
                           n_1116, QN => n1138);
   KEY_EXPAN0_reg_44_31_inst : FD1 port map( D => n6618, CP => CLK_I, Q => 
                           n_1117, QN => n67);
   KEY_EXPAN0_reg_43_31_inst : FD1 port map( D => n6617, CP => CLK_I, Q => 
                           n_1118, QN => n1137);
   KEY_EXPAN0_reg_42_31_inst : FD1 port map( D => n6616, CP => CLK_I, Q => 
                           n_1119, QN => n66);
   KEY_EXPAN0_reg_41_31_inst : FD1 port map( D => n6615, CP => CLK_I, Q => 
                           n_1120, QN => n1136);
   KEY_EXPAN0_reg_40_31_inst : FD1 port map( D => n6614, CP => CLK_I, Q => 
                           n_1121, QN => n65);
   KEY_EXPAN0_reg_39_31_inst : FD1 port map( D => n6613, CP => CLK_I, Q => 
                           n_1122, QN => n1143);
   KEY_EXPAN0_reg_38_31_inst : FD1 port map( D => n6612, CP => CLK_I, Q => 
                           n_1123, QN => n72);
   KEY_EXPAN0_reg_37_31_inst : FD1 port map( D => n6611, CP => CLK_I, Q => 
                           n_1124, QN => n1142);
   KEY_EXPAN0_reg_36_31_inst : FD1 port map( D => n6610, CP => CLK_I, Q => 
                           n_1125, QN => n71);
   KEY_EXPAN0_reg_35_31_inst : FD1 port map( D => n6609, CP => CLK_I, Q => 
                           n_1126, QN => n1141);
   KEY_EXPAN0_reg_34_31_inst : FD1 port map( D => n6608, CP => CLK_I, Q => 
                           n_1127, QN => n70);
   KEY_EXPAN0_reg_33_31_inst : FD1 port map( D => n6607, CP => CLK_I, Q => 
                           n_1128, QN => n1140);
   KEY_EXPAN0_reg_32_31_inst : FD1 port map( D => n6606, CP => CLK_I, Q => 
                           n_1129, QN => n69);
   KEY_EXPAN0_reg_31_31_inst : FD1 port map( D => n6605, CP => CLK_I, Q => 
                           n_1130, QN => n1115);
   KEY_EXPAN0_reg_30_31_inst : FD1 port map( D => n6604, CP => CLK_I, Q => 
                           n_1131, QN => n44);
   KEY_EXPAN0_reg_29_31_inst : FD1 port map( D => n6603, CP => CLK_I, Q => 
                           n_1132, QN => n1114);
   KEY_EXPAN0_reg_28_31_inst : FD1 port map( D => n6602, CP => CLK_I, Q => 
                           n_1133, QN => n43);
   KEY_EXPAN0_reg_27_31_inst : FD1 port map( D => n6601, CP => CLK_I, Q => 
                           n_1134, QN => n1113);
   KEY_EXPAN0_reg_26_31_inst : FD1 port map( D => n6600, CP => CLK_I, Q => 
                           n_1135, QN => n42);
   KEY_EXPAN0_reg_25_31_inst : FD1 port map( D => n6599, CP => CLK_I, Q => 
                           n_1136, QN => n1112);
   KEY_EXPAN0_reg_24_31_inst : FD1 port map( D => n6598, CP => CLK_I, Q => 
                           n_1137, QN => n41);
   KEY_EXPAN0_reg_23_31_inst : FD1 port map( D => n6597, CP => CLK_I, Q => 
                           n_1138, QN => n1119);
   KEY_EXPAN0_reg_22_31_inst : FD1 port map( D => n6596, CP => CLK_I, Q => 
                           n_1139, QN => n48);
   KEY_EXPAN0_reg_21_31_inst : FD1 port map( D => n6595, CP => CLK_I, Q => 
                           n_1140, QN => n1118);
   KEY_EXPAN0_reg_20_31_inst : FD1 port map( D => n6594, CP => CLK_I, Q => 
                           n_1141, QN => n47);
   KEY_EXPAN0_reg_19_31_inst : FD1 port map( D => n6593, CP => CLK_I, Q => 
                           n_1142, QN => n1117);
   KEY_EXPAN0_reg_18_31_inst : FD1 port map( D => n6592, CP => CLK_I, Q => 
                           n_1143, QN => n46);
   KEY_EXPAN0_reg_17_31_inst : FD1 port map( D => n6591, CP => CLK_I, Q => 
                           n_1144, QN => n1116);
   KEY_EXPAN0_reg_16_31_inst : FD1 port map( D => n6590, CP => CLK_I, Q => 
                           n_1145, QN => n45);
   KEY_EXPAN0_reg_15_31_inst : FD1 port map( D => n6589, CP => CLK_I, Q => 
                           n_1146, QN => n1123);
   KEY_EXPAN0_reg_14_31_inst : FD1 port map( D => n6588, CP => CLK_I, Q => 
                           n_1147, QN => n52);
   KEY_EXPAN0_reg_13_31_inst : FD1 port map( D => n6587, CP => CLK_I, Q => 
                           n_1148, QN => n1122);
   KEY_EXPAN0_reg_12_31_inst : FD1 port map( D => n6586, CP => CLK_I, Q => 
                           n_1149, QN => n51);
   KEY_EXPAN0_reg_11_31_inst : FD1 port map( D => n6585, CP => CLK_I, Q => 
                           n_1150, QN => n1121);
   KEY_EXPAN0_reg_10_31_inst : FD1 port map( D => n6584, CP => CLK_I, Q => 
                           n_1151, QN => n50);
   KEY_EXPAN0_reg_9_31_inst : FD1 port map( D => n6583, CP => CLK_I, Q => 
                           n_1152, QN => n1120);
   KEY_EXPAN0_reg_8_31_inst : FD1 port map( D => n6582, CP => CLK_I, Q => 
                           n_1153, QN => n49);
   KEY_EXPAN0_reg_7_31_inst : FD1 port map( D => n6581, CP => CLK_I, Q => 
                           n_1154, QN => n1127);
   KEY_EXPAN0_reg_6_31_inst : FD1 port map( D => n6580, CP => CLK_I, Q => 
                           n_1155, QN => n56);
   KEY_EXPAN0_reg_5_31_inst : FD1 port map( D => n6579, CP => CLK_I, Q => 
                           n_1156, QN => n1126);
   KEY_EXPAN0_reg_4_31_inst : FD1 port map( D => n6578, CP => CLK_I, Q => 
                           n_1157, QN => n55);
   KEY_EXPAN0_reg_3_31_inst : FD1 port map( D => n6577, CP => CLK_I, Q => 
                           n_1158, QN => n1125);
   KEY_EXPAN0_reg_2_31_inst : FD1 port map( D => n6576, CP => CLK_I, Q => 
                           n_1159, QN => n54);
   KEY_EXPAN0_reg_1_31_inst : FD1 port map( D => n6575, CP => CLK_I, Q => 
                           n_1160, QN => n1124);
   KEY_EXPAN0_reg_0_31_inst : FD1 port map( D => n6574, CP => CLK_I, Q => 
                           n_1161, QN => n53);
   v_KEY_COL_OUT0_reg_31_inst : FD1 port map( D => n4579, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_31_port, QN => n1050);
   v_TEMP_VECTOR_reg_23_inst : FD1 port map( D => n6672, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_23_port, QN => n_1162);
   KEY_EXPAN0_reg_63_23_inst : FD1 port map( D => n6125, CP => CLK_I, Q => 
                           n_1163, QN => n1163);
   KEY_EXPAN0_reg_62_23_inst : FD1 port map( D => n6124, CP => CLK_I, Q => 
                           n_1164, QN => n92);
   KEY_EXPAN0_reg_61_23_inst : FD1 port map( D => n6123, CP => CLK_I, Q => 
                           n_1165, QN => n1162);
   KEY_EXPAN0_reg_60_23_inst : FD1 port map( D => n6122, CP => CLK_I, Q => 
                           n_1166, QN => n91);
   KEY_EXPAN0_reg_59_23_inst : FD1 port map( D => n6121, CP => CLK_I, Q => 
                           n_1167, QN => n1161);
   KEY_EXPAN0_reg_58_23_inst : FD1 port map( D => n6120, CP => CLK_I, Q => 
                           n_1168, QN => n90);
   KEY_EXPAN0_reg_57_23_inst : FD1 port map( D => n6119, CP => CLK_I, Q => 
                           n_1169, QN => n1160);
   KEY_EXPAN0_reg_56_23_inst : FD1 port map( D => n6118, CP => CLK_I, Q => 
                           n_1170, QN => n89);
   KEY_EXPAN0_reg_55_23_inst : FD1 port map( D => n6117, CP => CLK_I, Q => 
                           n_1171, QN => n1167);
   KEY_EXPAN0_reg_54_23_inst : FD1 port map( D => n6116, CP => CLK_I, Q => 
                           n_1172, QN => n96);
   KEY_EXPAN0_reg_53_23_inst : FD1 port map( D => n6115, CP => CLK_I, Q => 
                           n_1173, QN => n1166);
   KEY_EXPAN0_reg_52_23_inst : FD1 port map( D => n6114, CP => CLK_I, Q => 
                           n_1174, QN => n95);
   KEY_EXPAN0_reg_51_23_inst : FD1 port map( D => n6113, CP => CLK_I, Q => 
                           n_1175, QN => n1165);
   KEY_EXPAN0_reg_50_23_inst : FD1 port map( D => n6112, CP => CLK_I, Q => 
                           n_1176, QN => n94);
   KEY_EXPAN0_reg_49_23_inst : FD1 port map( D => n6111, CP => CLK_I, Q => 
                           n_1177, QN => n1164);
   KEY_EXPAN0_reg_48_23_inst : FD1 port map( D => n6110, CP => CLK_I, Q => 
                           n_1178, QN => n93);
   KEY_EXPAN0_reg_47_23_inst : FD1 port map( D => n6109, CP => CLK_I, Q => 
                           n_1179, QN => n1171);
   KEY_EXPAN0_reg_46_23_inst : FD1 port map( D => n6108, CP => CLK_I, Q => 
                           n_1180, QN => n100);
   KEY_EXPAN0_reg_45_23_inst : FD1 port map( D => n6107, CP => CLK_I, Q => 
                           n_1181, QN => n1170);
   KEY_EXPAN0_reg_44_23_inst : FD1 port map( D => n6106, CP => CLK_I, Q => 
                           n_1182, QN => n99);
   KEY_EXPAN0_reg_43_23_inst : FD1 port map( D => n6105, CP => CLK_I, Q => 
                           n_1183, QN => n1169);
   KEY_EXPAN0_reg_42_23_inst : FD1 port map( D => n6104, CP => CLK_I, Q => 
                           n_1184, QN => n98);
   KEY_EXPAN0_reg_41_23_inst : FD1 port map( D => n6103, CP => CLK_I, Q => 
                           n_1185, QN => n1168);
   KEY_EXPAN0_reg_40_23_inst : FD1 port map( D => n6102, CP => CLK_I, Q => 
                           n_1186, QN => n97);
   KEY_EXPAN0_reg_39_23_inst : FD1 port map( D => n6101, CP => CLK_I, Q => 
                           n_1187, QN => n1175);
   KEY_EXPAN0_reg_38_23_inst : FD1 port map( D => n6100, CP => CLK_I, Q => 
                           n_1188, QN => n104);
   KEY_EXPAN0_reg_37_23_inst : FD1 port map( D => n6099, CP => CLK_I, Q => 
                           n_1189, QN => n1174);
   KEY_EXPAN0_reg_36_23_inst : FD1 port map( D => n6098, CP => CLK_I, Q => 
                           n_1190, QN => n103);
   KEY_EXPAN0_reg_35_23_inst : FD1 port map( D => n6097, CP => CLK_I, Q => 
                           n_1191, QN => n1173);
   KEY_EXPAN0_reg_34_23_inst : FD1 port map( D => n6096, CP => CLK_I, Q => 
                           n_1192, QN => n102);
   KEY_EXPAN0_reg_33_23_inst : FD1 port map( D => n6095, CP => CLK_I, Q => 
                           n_1193, QN => n1172);
   KEY_EXPAN0_reg_32_23_inst : FD1 port map( D => n6094, CP => CLK_I, Q => 
                           n_1194, QN => n101);
   KEY_EXPAN0_reg_31_23_inst : FD1 port map( D => n6093, CP => CLK_I, Q => 
                           n_1195, QN => n1147);
   KEY_EXPAN0_reg_30_23_inst : FD1 port map( D => n6092, CP => CLK_I, Q => 
                           n_1196, QN => n76);
   KEY_EXPAN0_reg_29_23_inst : FD1 port map( D => n6091, CP => CLK_I, Q => 
                           n_1197, QN => n1146);
   KEY_EXPAN0_reg_28_23_inst : FD1 port map( D => n6090, CP => CLK_I, Q => 
                           n_1198, QN => n75);
   KEY_EXPAN0_reg_27_23_inst : FD1 port map( D => n6089, CP => CLK_I, Q => 
                           n_1199, QN => n1145);
   KEY_EXPAN0_reg_26_23_inst : FD1 port map( D => n6088, CP => CLK_I, Q => 
                           n_1200, QN => n74);
   KEY_EXPAN0_reg_25_23_inst : FD1 port map( D => n6087, CP => CLK_I, Q => 
                           n_1201, QN => n1144);
   KEY_EXPAN0_reg_24_23_inst : FD1 port map( D => n6086, CP => CLK_I, Q => 
                           n_1202, QN => n73);
   KEY_EXPAN0_reg_23_23_inst : FD1 port map( D => n6085, CP => CLK_I, Q => 
                           n_1203, QN => n1151);
   KEY_EXPAN0_reg_22_23_inst : FD1 port map( D => n6084, CP => CLK_I, Q => 
                           n_1204, QN => n80);
   KEY_EXPAN0_reg_21_23_inst : FD1 port map( D => n6083, CP => CLK_I, Q => 
                           n_1205, QN => n1150);
   KEY_EXPAN0_reg_20_23_inst : FD1 port map( D => n6082, CP => CLK_I, Q => 
                           n_1206, QN => n79);
   KEY_EXPAN0_reg_19_23_inst : FD1 port map( D => n6081, CP => CLK_I, Q => 
                           n_1207, QN => n1149);
   KEY_EXPAN0_reg_18_23_inst : FD1 port map( D => n6080, CP => CLK_I, Q => 
                           n_1208, QN => n78);
   KEY_EXPAN0_reg_17_23_inst : FD1 port map( D => n6079, CP => CLK_I, Q => 
                           n_1209, QN => n1148);
   KEY_EXPAN0_reg_16_23_inst : FD1 port map( D => n6078, CP => CLK_I, Q => 
                           n_1210, QN => n77);
   KEY_EXPAN0_reg_15_23_inst : FD1 port map( D => n6077, CP => CLK_I, Q => 
                           n_1211, QN => n1155);
   KEY_EXPAN0_reg_14_23_inst : FD1 port map( D => n6076, CP => CLK_I, Q => 
                           n_1212, QN => n84);
   KEY_EXPAN0_reg_13_23_inst : FD1 port map( D => n6075, CP => CLK_I, Q => 
                           n_1213, QN => n1154);
   KEY_EXPAN0_reg_12_23_inst : FD1 port map( D => n6074, CP => CLK_I, Q => 
                           n_1214, QN => n83);
   KEY_EXPAN0_reg_11_23_inst : FD1 port map( D => n6073, CP => CLK_I, Q => 
                           n_1215, QN => n1153);
   KEY_EXPAN0_reg_10_23_inst : FD1 port map( D => n6072, CP => CLK_I, Q => 
                           n_1216, QN => n82);
   KEY_EXPAN0_reg_9_23_inst : FD1 port map( D => n6071, CP => CLK_I, Q => 
                           n_1217, QN => n1152);
   KEY_EXPAN0_reg_8_23_inst : FD1 port map( D => n6070, CP => CLK_I, Q => 
                           n_1218, QN => n81);
   KEY_EXPAN0_reg_7_23_inst : FD1 port map( D => n6069, CP => CLK_I, Q => 
                           n_1219, QN => n1159);
   KEY_EXPAN0_reg_6_23_inst : FD1 port map( D => n6068, CP => CLK_I, Q => 
                           n_1220, QN => n88);
   KEY_EXPAN0_reg_5_23_inst : FD1 port map( D => n6067, CP => CLK_I, Q => 
                           n_1221, QN => n1158);
   KEY_EXPAN0_reg_4_23_inst : FD1 port map( D => n6066, CP => CLK_I, Q => 
                           n_1222, QN => n87);
   KEY_EXPAN0_reg_3_23_inst : FD1 port map( D => n6065, CP => CLK_I, Q => 
                           n_1223, QN => n1157);
   KEY_EXPAN0_reg_2_23_inst : FD1 port map( D => n6064, CP => CLK_I, Q => 
                           n_1224, QN => n86);
   KEY_EXPAN0_reg_1_23_inst : FD1 port map( D => n6063, CP => CLK_I, Q => 
                           n_1225, QN => n1156);
   KEY_EXPAN0_reg_0_23_inst : FD1 port map( D => n6062, CP => CLK_I, Q => 
                           n_1226, QN => n85);
   v_KEY_COL_OUT0_reg_23_inst : FD1 port map( D => n4578, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_23_port, QN => n1059);
   v_TEMP_VECTOR_reg_15_inst : FD1 port map( D => n6680, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_15_port, QN => n_1227);
   KEY_EXPAN0_reg_63_15_inst : FD1 port map( D => n5613, CP => CLK_I, Q => 
                           n_1228, QN => n1195);
   KEY_EXPAN0_reg_62_15_inst : FD1 port map( D => n5612, CP => CLK_I, Q => 
                           n_1229, QN => n124);
   KEY_EXPAN0_reg_61_15_inst : FD1 port map( D => n5611, CP => CLK_I, Q => 
                           n_1230, QN => n1194);
   KEY_EXPAN0_reg_60_15_inst : FD1 port map( D => n5610, CP => CLK_I, Q => 
                           n_1231, QN => n123);
   KEY_EXPAN0_reg_59_15_inst : FD1 port map( D => n5609, CP => CLK_I, Q => 
                           n_1232, QN => n1193);
   KEY_EXPAN0_reg_58_15_inst : FD1 port map( D => n5608, CP => CLK_I, Q => 
                           n_1233, QN => n122);
   KEY_EXPAN0_reg_57_15_inst : FD1 port map( D => n5607, CP => CLK_I, Q => 
                           n_1234, QN => n1192);
   KEY_EXPAN0_reg_56_15_inst : FD1 port map( D => n5606, CP => CLK_I, Q => 
                           n_1235, QN => n121);
   KEY_EXPAN0_reg_55_15_inst : FD1 port map( D => n5605, CP => CLK_I, Q => 
                           n_1236, QN => n1199);
   KEY_EXPAN0_reg_54_15_inst : FD1 port map( D => n5604, CP => CLK_I, Q => 
                           n_1237, QN => n128);
   KEY_EXPAN0_reg_53_15_inst : FD1 port map( D => n5603, CP => CLK_I, Q => 
                           n_1238, QN => n1198);
   KEY_EXPAN0_reg_52_15_inst : FD1 port map( D => n5602, CP => CLK_I, Q => 
                           n_1239, QN => n127);
   KEY_EXPAN0_reg_51_15_inst : FD1 port map( D => n5601, CP => CLK_I, Q => 
                           n_1240, QN => n1197);
   KEY_EXPAN0_reg_50_15_inst : FD1 port map( D => n5600, CP => CLK_I, Q => 
                           n_1241, QN => n126);
   KEY_EXPAN0_reg_49_15_inst : FD1 port map( D => n5599, CP => CLK_I, Q => 
                           n_1242, QN => n1196);
   KEY_EXPAN0_reg_48_15_inst : FD1 port map( D => n5598, CP => CLK_I, Q => 
                           n_1243, QN => n125);
   KEY_EXPAN0_reg_47_15_inst : FD1 port map( D => n5597, CP => CLK_I, Q => 
                           n_1244, QN => n1203);
   KEY_EXPAN0_reg_46_15_inst : FD1 port map( D => n5596, CP => CLK_I, Q => 
                           n_1245, QN => n132);
   KEY_EXPAN0_reg_45_15_inst : FD1 port map( D => n5595, CP => CLK_I, Q => 
                           n_1246, QN => n1202);
   KEY_EXPAN0_reg_44_15_inst : FD1 port map( D => n5594, CP => CLK_I, Q => 
                           n_1247, QN => n131);
   KEY_EXPAN0_reg_43_15_inst : FD1 port map( D => n5593, CP => CLK_I, Q => 
                           n_1248, QN => n1201);
   KEY_EXPAN0_reg_42_15_inst : FD1 port map( D => n5592, CP => CLK_I, Q => 
                           n_1249, QN => n130);
   KEY_EXPAN0_reg_41_15_inst : FD1 port map( D => n5591, CP => CLK_I, Q => 
                           n_1250, QN => n1200);
   KEY_EXPAN0_reg_40_15_inst : FD1 port map( D => n5590, CP => CLK_I, Q => 
                           n_1251, QN => n129);
   KEY_EXPAN0_reg_39_15_inst : FD1 port map( D => n5589, CP => CLK_I, Q => 
                           n_1252, QN => n1207);
   KEY_EXPAN0_reg_38_15_inst : FD1 port map( D => n5588, CP => CLK_I, Q => 
                           n_1253, QN => n136);
   KEY_EXPAN0_reg_37_15_inst : FD1 port map( D => n5587, CP => CLK_I, Q => 
                           n_1254, QN => n1206);
   KEY_EXPAN0_reg_36_15_inst : FD1 port map( D => n5586, CP => CLK_I, Q => 
                           n_1255, QN => n135);
   KEY_EXPAN0_reg_35_15_inst : FD1 port map( D => n5585, CP => CLK_I, Q => 
                           n_1256, QN => n1205);
   KEY_EXPAN0_reg_34_15_inst : FD1 port map( D => n5584, CP => CLK_I, Q => 
                           n_1257, QN => n134);
   KEY_EXPAN0_reg_33_15_inst : FD1 port map( D => n5583, CP => CLK_I, Q => 
                           n_1258, QN => n1204);
   KEY_EXPAN0_reg_32_15_inst : FD1 port map( D => n5582, CP => CLK_I, Q => 
                           n_1259, QN => n133);
   KEY_EXPAN0_reg_31_15_inst : FD1 port map( D => n5581, CP => CLK_I, Q => 
                           n_1260, QN => n1179);
   KEY_EXPAN0_reg_30_15_inst : FD1 port map( D => n5580, CP => CLK_I, Q => 
                           n_1261, QN => n108);
   KEY_EXPAN0_reg_29_15_inst : FD1 port map( D => n5579, CP => CLK_I, Q => 
                           n_1262, QN => n1178);
   KEY_EXPAN0_reg_28_15_inst : FD1 port map( D => n5578, CP => CLK_I, Q => 
                           n_1263, QN => n107);
   KEY_EXPAN0_reg_27_15_inst : FD1 port map( D => n5577, CP => CLK_I, Q => 
                           n_1264, QN => n1177);
   KEY_EXPAN0_reg_26_15_inst : FD1 port map( D => n5576, CP => CLK_I, Q => 
                           n_1265, QN => n106);
   KEY_EXPAN0_reg_25_15_inst : FD1 port map( D => n5575, CP => CLK_I, Q => 
                           n_1266, QN => n1176);
   KEY_EXPAN0_reg_24_15_inst : FD1 port map( D => n5574, CP => CLK_I, Q => 
                           n_1267, QN => n105);
   KEY_EXPAN0_reg_23_15_inst : FD1 port map( D => n5573, CP => CLK_I, Q => 
                           n_1268, QN => n1183);
   KEY_EXPAN0_reg_22_15_inst : FD1 port map( D => n5572, CP => CLK_I, Q => 
                           n_1269, QN => n112);
   KEY_EXPAN0_reg_21_15_inst : FD1 port map( D => n5571, CP => CLK_I, Q => 
                           n_1270, QN => n1182);
   KEY_EXPAN0_reg_20_15_inst : FD1 port map( D => n5570, CP => CLK_I, Q => 
                           n_1271, QN => n111);
   KEY_EXPAN0_reg_19_15_inst : FD1 port map( D => n5569, CP => CLK_I, Q => 
                           n_1272, QN => n1181);
   KEY_EXPAN0_reg_18_15_inst : FD1 port map( D => n5568, CP => CLK_I, Q => 
                           n_1273, QN => n110);
   KEY_EXPAN0_reg_17_15_inst : FD1 port map( D => n5567, CP => CLK_I, Q => 
                           n_1274, QN => n1180);
   KEY_EXPAN0_reg_16_15_inst : FD1 port map( D => n5566, CP => CLK_I, Q => 
                           n_1275, QN => n109);
   KEY_EXPAN0_reg_15_15_inst : FD1 port map( D => n5565, CP => CLK_I, Q => 
                           n_1276, QN => n1187);
   KEY_EXPAN0_reg_14_15_inst : FD1 port map( D => n5564, CP => CLK_I, Q => 
                           n_1277, QN => n116);
   KEY_EXPAN0_reg_13_15_inst : FD1 port map( D => n5563, CP => CLK_I, Q => 
                           n_1278, QN => n1186);
   KEY_EXPAN0_reg_12_15_inst : FD1 port map( D => n5562, CP => CLK_I, Q => 
                           n_1279, QN => n115);
   KEY_EXPAN0_reg_11_15_inst : FD1 port map( D => n5561, CP => CLK_I, Q => 
                           n_1280, QN => n1185);
   KEY_EXPAN0_reg_10_15_inst : FD1 port map( D => n5560, CP => CLK_I, Q => 
                           n_1281, QN => n114);
   KEY_EXPAN0_reg_9_15_inst : FD1 port map( D => n5559, CP => CLK_I, Q => 
                           n_1282, QN => n1184);
   KEY_EXPAN0_reg_8_15_inst : FD1 port map( D => n5558, CP => CLK_I, Q => 
                           n_1283, QN => n113);
   KEY_EXPAN0_reg_7_15_inst : FD1 port map( D => n5557, CP => CLK_I, Q => 
                           n_1284, QN => n1191);
   KEY_EXPAN0_reg_6_15_inst : FD1 port map( D => n5556, CP => CLK_I, Q => 
                           n_1285, QN => n120);
   KEY_EXPAN0_reg_5_15_inst : FD1 port map( D => n5555, CP => CLK_I, Q => 
                           n_1286, QN => n1190);
   KEY_EXPAN0_reg_4_15_inst : FD1 port map( D => n5554, CP => CLK_I, Q => 
                           n_1287, QN => n119);
   KEY_EXPAN0_reg_3_15_inst : FD1 port map( D => n5553, CP => CLK_I, Q => 
                           n_1288, QN => n1189);
   KEY_EXPAN0_reg_2_15_inst : FD1 port map( D => n5552, CP => CLK_I, Q => 
                           n_1289, QN => n118);
   KEY_EXPAN0_reg_1_15_inst : FD1 port map( D => n5551, CP => CLK_I, Q => 
                           n_1290, QN => n1188);
   KEY_EXPAN0_reg_0_15_inst : FD1 port map( D => n5550, CP => CLK_I, Q => 
                           n_1291, QN => n117);
   v_KEY_COL_OUT0_reg_15_inst : FD1 port map( D => n4577, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_15_port, QN => n1068);
   v_TEMP_VECTOR_reg_6_inst : FD1 port map( D => n6689, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_6_port, QN => n_1292);
   KEY_EXPAN0_reg_63_6_inst : FD1 port map( D => n5037, CP => CLK_I, Q => 
                           n_1293, QN => n1227);
   KEY_EXPAN0_reg_62_6_inst : FD1 port map( D => n5036, CP => CLK_I, Q => 
                           n_1294, QN => n156);
   KEY_EXPAN0_reg_61_6_inst : FD1 port map( D => n5035, CP => CLK_I, Q => 
                           n_1295, QN => n1226);
   KEY_EXPAN0_reg_60_6_inst : FD1 port map( D => n5034, CP => CLK_I, Q => 
                           n_1296, QN => n155);
   KEY_EXPAN0_reg_59_6_inst : FD1 port map( D => n5033, CP => CLK_I, Q => 
                           n_1297, QN => n1225);
   KEY_EXPAN0_reg_58_6_inst : FD1 port map( D => n5032, CP => CLK_I, Q => 
                           n_1298, QN => n154);
   KEY_EXPAN0_reg_57_6_inst : FD1 port map( D => n5031, CP => CLK_I, Q => 
                           n_1299, QN => n1224);
   KEY_EXPAN0_reg_56_6_inst : FD1 port map( D => n5030, CP => CLK_I, Q => 
                           n_1300, QN => n153);
   KEY_EXPAN0_reg_55_6_inst : FD1 port map( D => n5029, CP => CLK_I, Q => 
                           n_1301, QN => n1231);
   KEY_EXPAN0_reg_54_6_inst : FD1 port map( D => n5028, CP => CLK_I, Q => 
                           n_1302, QN => n160);
   KEY_EXPAN0_reg_53_6_inst : FD1 port map( D => n5027, CP => CLK_I, Q => 
                           n_1303, QN => n1230);
   KEY_EXPAN0_reg_52_6_inst : FD1 port map( D => n5026, CP => CLK_I, Q => 
                           n_1304, QN => n159);
   KEY_EXPAN0_reg_51_6_inst : FD1 port map( D => n5025, CP => CLK_I, Q => 
                           n_1305, QN => n1229);
   KEY_EXPAN0_reg_50_6_inst : FD1 port map( D => n5024, CP => CLK_I, Q => 
                           n_1306, QN => n158);
   KEY_EXPAN0_reg_49_6_inst : FD1 port map( D => n5023, CP => CLK_I, Q => 
                           n_1307, QN => n1228);
   KEY_EXPAN0_reg_48_6_inst : FD1 port map( D => n5022, CP => CLK_I, Q => 
                           n_1308, QN => n157);
   KEY_EXPAN0_reg_47_6_inst : FD1 port map( D => n5021, CP => CLK_I, Q => 
                           n_1309, QN => n1235);
   KEY_EXPAN0_reg_46_6_inst : FD1 port map( D => n5020, CP => CLK_I, Q => 
                           n_1310, QN => n164);
   KEY_EXPAN0_reg_45_6_inst : FD1 port map( D => n5019, CP => CLK_I, Q => 
                           n_1311, QN => n1234);
   KEY_EXPAN0_reg_44_6_inst : FD1 port map( D => n5018, CP => CLK_I, Q => 
                           n_1312, QN => n163);
   KEY_EXPAN0_reg_43_6_inst : FD1 port map( D => n5017, CP => CLK_I, Q => 
                           n_1313, QN => n1233);
   KEY_EXPAN0_reg_42_6_inst : FD1 port map( D => n5016, CP => CLK_I, Q => 
                           n_1314, QN => n162);
   KEY_EXPAN0_reg_41_6_inst : FD1 port map( D => n5015, CP => CLK_I, Q => 
                           n_1315, QN => n1232);
   KEY_EXPAN0_reg_40_6_inst : FD1 port map( D => n5014, CP => CLK_I, Q => 
                           n_1316, QN => n161);
   KEY_EXPAN0_reg_39_6_inst : FD1 port map( D => n5013, CP => CLK_I, Q => 
                           n_1317, QN => n1239);
   KEY_EXPAN0_reg_38_6_inst : FD1 port map( D => n5012, CP => CLK_I, Q => 
                           n_1318, QN => n168);
   KEY_EXPAN0_reg_37_6_inst : FD1 port map( D => n5011, CP => CLK_I, Q => 
                           n_1319, QN => n1238);
   KEY_EXPAN0_reg_36_6_inst : FD1 port map( D => n5010, CP => CLK_I, Q => 
                           n_1320, QN => n167);
   KEY_EXPAN0_reg_35_6_inst : FD1 port map( D => n5009, CP => CLK_I, Q => 
                           n_1321, QN => n1237);
   KEY_EXPAN0_reg_34_6_inst : FD1 port map( D => n5008, CP => CLK_I, Q => 
                           n_1322, QN => n166);
   KEY_EXPAN0_reg_33_6_inst : FD1 port map( D => n5007, CP => CLK_I, Q => 
                           n_1323, QN => n1236);
   KEY_EXPAN0_reg_32_6_inst : FD1 port map( D => n5006, CP => CLK_I, Q => 
                           n_1324, QN => n165);
   KEY_EXPAN0_reg_31_6_inst : FD1 port map( D => n5005, CP => CLK_I, Q => 
                           n_1325, QN => n1211);
   KEY_EXPAN0_reg_30_6_inst : FD1 port map( D => n5004, CP => CLK_I, Q => 
                           n_1326, QN => n140);
   KEY_EXPAN0_reg_29_6_inst : FD1 port map( D => n5003, CP => CLK_I, Q => 
                           n_1327, QN => n1210);
   KEY_EXPAN0_reg_28_6_inst : FD1 port map( D => n5002, CP => CLK_I, Q => 
                           n_1328, QN => n139);
   KEY_EXPAN0_reg_27_6_inst : FD1 port map( D => n5001, CP => CLK_I, Q => 
                           n_1329, QN => n1209);
   KEY_EXPAN0_reg_26_6_inst : FD1 port map( D => n5000, CP => CLK_I, Q => 
                           n_1330, QN => n138);
   KEY_EXPAN0_reg_25_6_inst : FD1 port map( D => n4999, CP => CLK_I, Q => 
                           n_1331, QN => n1208);
   KEY_EXPAN0_reg_24_6_inst : FD1 port map( D => n4998, CP => CLK_I, Q => 
                           n_1332, QN => n137);
   KEY_EXPAN0_reg_23_6_inst : FD1 port map( D => n4997, CP => CLK_I, Q => 
                           n_1333, QN => n1215);
   KEY_EXPAN0_reg_22_6_inst : FD1 port map( D => n4996, CP => CLK_I, Q => 
                           n_1334, QN => n144);
   KEY_EXPAN0_reg_21_6_inst : FD1 port map( D => n4995, CP => CLK_I, Q => 
                           n_1335, QN => n1214);
   KEY_EXPAN0_reg_20_6_inst : FD1 port map( D => n4994, CP => CLK_I, Q => 
                           n_1336, QN => n143);
   KEY_EXPAN0_reg_19_6_inst : FD1 port map( D => n4993, CP => CLK_I, Q => 
                           n_1337, QN => n1213);
   KEY_EXPAN0_reg_18_6_inst : FD1 port map( D => n4992, CP => CLK_I, Q => 
                           n_1338, QN => n142);
   KEY_EXPAN0_reg_17_6_inst : FD1 port map( D => n4991, CP => CLK_I, Q => 
                           n_1339, QN => n1212);
   KEY_EXPAN0_reg_16_6_inst : FD1 port map( D => n4990, CP => CLK_I, Q => 
                           n_1340, QN => n141);
   KEY_EXPAN0_reg_15_6_inst : FD1 port map( D => n4989, CP => CLK_I, Q => 
                           n_1341, QN => n1219);
   KEY_EXPAN0_reg_14_6_inst : FD1 port map( D => n4988, CP => CLK_I, Q => 
                           n_1342, QN => n148);
   KEY_EXPAN0_reg_13_6_inst : FD1 port map( D => n4987, CP => CLK_I, Q => 
                           n_1343, QN => n1218);
   KEY_EXPAN0_reg_12_6_inst : FD1 port map( D => n4986, CP => CLK_I, Q => 
                           n_1344, QN => n147);
   KEY_EXPAN0_reg_11_6_inst : FD1 port map( D => n4985, CP => CLK_I, Q => 
                           n_1345, QN => n1217);
   KEY_EXPAN0_reg_10_6_inst : FD1 port map( D => n4984, CP => CLK_I, Q => 
                           n_1346, QN => n146);
   KEY_EXPAN0_reg_9_6_inst : FD1 port map( D => n4983, CP => CLK_I, Q => n_1347
                           , QN => n1216);
   KEY_EXPAN0_reg_8_6_inst : FD1 port map( D => n4982, CP => CLK_I, Q => n_1348
                           , QN => n145);
   KEY_EXPAN0_reg_7_6_inst : FD1 port map( D => n4981, CP => CLK_I, Q => n_1349
                           , QN => n1223);
   KEY_EXPAN0_reg_6_6_inst : FD1 port map( D => n4980, CP => CLK_I, Q => n_1350
                           , QN => n152);
   KEY_EXPAN0_reg_5_6_inst : FD1 port map( D => n4979, CP => CLK_I, Q => n_1351
                           , QN => n1222);
   KEY_EXPAN0_reg_4_6_inst : FD1 port map( D => n4978, CP => CLK_I, Q => n_1352
                           , QN => n151);
   KEY_EXPAN0_reg_3_6_inst : FD1 port map( D => n4977, CP => CLK_I, Q => n_1353
                           , QN => n1221);
   KEY_EXPAN0_reg_2_6_inst : FD1 port map( D => n4976, CP => CLK_I, Q => n_1354
                           , QN => n150);
   KEY_EXPAN0_reg_1_6_inst : FD1 port map( D => n4975, CP => CLK_I, Q => n_1355
                           , QN => n1220);
   KEY_EXPAN0_reg_0_6_inst : FD1 port map( D => n4974, CP => CLK_I, Q => n_1356
                           , QN => n149);
   v_KEY_COL_OUT0_reg_6_inst : FD1 port map( D => n4576, CP => CLK_I, Q => 
                           n2118, QN => n4457);
   v_TEMP_VECTOR_reg_30_inst : FD1 port map( D => n6665, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_30_port, QN => n_1357);
   KEY_EXPAN0_reg_63_30_inst : FD1 port map( D => n6573, CP => CLK_I, Q => 
                           n_1358, QN => n1259);
   KEY_EXPAN0_reg_62_30_inst : FD1 port map( D => n6572, CP => CLK_I, Q => 
                           n_1359, QN => n188);
   KEY_EXPAN0_reg_61_30_inst : FD1 port map( D => n6571, CP => CLK_I, Q => 
                           n_1360, QN => n1258);
   KEY_EXPAN0_reg_60_30_inst : FD1 port map( D => n6570, CP => CLK_I, Q => 
                           n_1361, QN => n187);
   KEY_EXPAN0_reg_59_30_inst : FD1 port map( D => n6569, CP => CLK_I, Q => 
                           n_1362, QN => n1257);
   KEY_EXPAN0_reg_58_30_inst : FD1 port map( D => n6568, CP => CLK_I, Q => 
                           n_1363, QN => n186);
   KEY_EXPAN0_reg_57_30_inst : FD1 port map( D => n6567, CP => CLK_I, Q => 
                           n_1364, QN => n1256);
   KEY_EXPAN0_reg_56_30_inst : FD1 port map( D => n6566, CP => CLK_I, Q => 
                           n_1365, QN => n185);
   KEY_EXPAN0_reg_55_30_inst : FD1 port map( D => n6565, CP => CLK_I, Q => 
                           n_1366, QN => n1263);
   KEY_EXPAN0_reg_54_30_inst : FD1 port map( D => n6564, CP => CLK_I, Q => 
                           n_1367, QN => n192);
   KEY_EXPAN0_reg_53_30_inst : FD1 port map( D => n6563, CP => CLK_I, Q => 
                           n_1368, QN => n1262);
   KEY_EXPAN0_reg_52_30_inst : FD1 port map( D => n6562, CP => CLK_I, Q => 
                           n_1369, QN => n191);
   KEY_EXPAN0_reg_51_30_inst : FD1 port map( D => n6561, CP => CLK_I, Q => 
                           n_1370, QN => n1261);
   KEY_EXPAN0_reg_50_30_inst : FD1 port map( D => n6560, CP => CLK_I, Q => 
                           n_1371, QN => n190);
   KEY_EXPAN0_reg_49_30_inst : FD1 port map( D => n6559, CP => CLK_I, Q => 
                           n_1372, QN => n1260);
   KEY_EXPAN0_reg_48_30_inst : FD1 port map( D => n6558, CP => CLK_I, Q => 
                           n_1373, QN => n189);
   KEY_EXPAN0_reg_47_30_inst : FD1 port map( D => n6557, CP => CLK_I, Q => 
                           n_1374, QN => n1267);
   KEY_EXPAN0_reg_46_30_inst : FD1 port map( D => n6556, CP => CLK_I, Q => 
                           n_1375, QN => n196);
   KEY_EXPAN0_reg_45_30_inst : FD1 port map( D => n6555, CP => CLK_I, Q => 
                           n_1376, QN => n1266);
   KEY_EXPAN0_reg_44_30_inst : FD1 port map( D => n6554, CP => CLK_I, Q => 
                           n_1377, QN => n195);
   KEY_EXPAN0_reg_43_30_inst : FD1 port map( D => n6553, CP => CLK_I, Q => 
                           n_1378, QN => n1265);
   KEY_EXPAN0_reg_42_30_inst : FD1 port map( D => n6552, CP => CLK_I, Q => 
                           n_1379, QN => n194);
   KEY_EXPAN0_reg_41_30_inst : FD1 port map( D => n6551, CP => CLK_I, Q => 
                           n_1380, QN => n1264);
   KEY_EXPAN0_reg_40_30_inst : FD1 port map( D => n6550, CP => CLK_I, Q => 
                           n_1381, QN => n193);
   KEY_EXPAN0_reg_39_30_inst : FD1 port map( D => n6549, CP => CLK_I, Q => 
                           n_1382, QN => n1271);
   KEY_EXPAN0_reg_38_30_inst : FD1 port map( D => n6548, CP => CLK_I, Q => 
                           n_1383, QN => n200);
   KEY_EXPAN0_reg_37_30_inst : FD1 port map( D => n6547, CP => CLK_I, Q => 
                           n_1384, QN => n1270);
   KEY_EXPAN0_reg_36_30_inst : FD1 port map( D => n6546, CP => CLK_I, Q => 
                           n_1385, QN => n199);
   KEY_EXPAN0_reg_35_30_inst : FD1 port map( D => n6545, CP => CLK_I, Q => 
                           n_1386, QN => n1269);
   KEY_EXPAN0_reg_34_30_inst : FD1 port map( D => n6544, CP => CLK_I, Q => 
                           n_1387, QN => n198);
   KEY_EXPAN0_reg_33_30_inst : FD1 port map( D => n6543, CP => CLK_I, Q => 
                           n_1388, QN => n1268);
   KEY_EXPAN0_reg_32_30_inst : FD1 port map( D => n6542, CP => CLK_I, Q => 
                           n_1389, QN => n197);
   KEY_EXPAN0_reg_31_30_inst : FD1 port map( D => n6541, CP => CLK_I, Q => 
                           n_1390, QN => n1243);
   KEY_EXPAN0_reg_30_30_inst : FD1 port map( D => n6540, CP => CLK_I, Q => 
                           n_1391, QN => n172);
   KEY_EXPAN0_reg_29_30_inst : FD1 port map( D => n6539, CP => CLK_I, Q => 
                           n_1392, QN => n1242);
   KEY_EXPAN0_reg_28_30_inst : FD1 port map( D => n6538, CP => CLK_I, Q => 
                           n_1393, QN => n171);
   KEY_EXPAN0_reg_27_30_inst : FD1 port map( D => n6537, CP => CLK_I, Q => 
                           n_1394, QN => n1241);
   KEY_EXPAN0_reg_26_30_inst : FD1 port map( D => n6536, CP => CLK_I, Q => 
                           n_1395, QN => n170);
   KEY_EXPAN0_reg_25_30_inst : FD1 port map( D => n6535, CP => CLK_I, Q => 
                           n_1396, QN => n1240);
   KEY_EXPAN0_reg_24_30_inst : FD1 port map( D => n6534, CP => CLK_I, Q => 
                           n_1397, QN => n169);
   KEY_EXPAN0_reg_23_30_inst : FD1 port map( D => n6533, CP => CLK_I, Q => 
                           n_1398, QN => n1247);
   KEY_EXPAN0_reg_22_30_inst : FD1 port map( D => n6532, CP => CLK_I, Q => 
                           n_1399, QN => n176);
   KEY_EXPAN0_reg_21_30_inst : FD1 port map( D => n6531, CP => CLK_I, Q => 
                           n_1400, QN => n1246);
   KEY_EXPAN0_reg_20_30_inst : FD1 port map( D => n6530, CP => CLK_I, Q => 
                           n_1401, QN => n175);
   KEY_EXPAN0_reg_19_30_inst : FD1 port map( D => n6529, CP => CLK_I, Q => 
                           n_1402, QN => n1245);
   KEY_EXPAN0_reg_18_30_inst : FD1 port map( D => n6528, CP => CLK_I, Q => 
                           n_1403, QN => n174);
   KEY_EXPAN0_reg_17_30_inst : FD1 port map( D => n6527, CP => CLK_I, Q => 
                           n_1404, QN => n1244);
   KEY_EXPAN0_reg_16_30_inst : FD1 port map( D => n6526, CP => CLK_I, Q => 
                           n_1405, QN => n173);
   KEY_EXPAN0_reg_15_30_inst : FD1 port map( D => n6525, CP => CLK_I, Q => 
                           n_1406, QN => n1251);
   KEY_EXPAN0_reg_14_30_inst : FD1 port map( D => n6524, CP => CLK_I, Q => 
                           n_1407, QN => n180);
   KEY_EXPAN0_reg_13_30_inst : FD1 port map( D => n6523, CP => CLK_I, Q => 
                           n_1408, QN => n1250);
   KEY_EXPAN0_reg_12_30_inst : FD1 port map( D => n6522, CP => CLK_I, Q => 
                           n_1409, QN => n179);
   KEY_EXPAN0_reg_11_30_inst : FD1 port map( D => n6521, CP => CLK_I, Q => 
                           n_1410, QN => n1249);
   KEY_EXPAN0_reg_10_30_inst : FD1 port map( D => n6520, CP => CLK_I, Q => 
                           n_1411, QN => n178);
   KEY_EXPAN0_reg_9_30_inst : FD1 port map( D => n6519, CP => CLK_I, Q => 
                           n_1412, QN => n1248);
   KEY_EXPAN0_reg_8_30_inst : FD1 port map( D => n6518, CP => CLK_I, Q => 
                           n_1413, QN => n177);
   KEY_EXPAN0_reg_7_30_inst : FD1 port map( D => n6517, CP => CLK_I, Q => 
                           n_1414, QN => n1255);
   KEY_EXPAN0_reg_6_30_inst : FD1 port map( D => n6516, CP => CLK_I, Q => 
                           n_1415, QN => n184);
   KEY_EXPAN0_reg_5_30_inst : FD1 port map( D => n6515, CP => CLK_I, Q => 
                           n_1416, QN => n1254);
   KEY_EXPAN0_reg_4_30_inst : FD1 port map( D => n6514, CP => CLK_I, Q => 
                           n_1417, QN => n183);
   KEY_EXPAN0_reg_3_30_inst : FD1 port map( D => n6513, CP => CLK_I, Q => 
                           n_1418, QN => n1253);
   KEY_EXPAN0_reg_2_30_inst : FD1 port map( D => n6512, CP => CLK_I, Q => 
                           n_1419, QN => n182);
   KEY_EXPAN0_reg_1_30_inst : FD1 port map( D => n6511, CP => CLK_I, Q => 
                           n_1420, QN => n1252);
   KEY_EXPAN0_reg_0_30_inst : FD1 port map( D => n6510, CP => CLK_I, Q => 
                           n_1421, QN => n181);
   v_KEY_COL_OUT0_reg_30_inst : FD1 port map( D => n4575, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_30_port, QN => n1051);
   v_TEMP_VECTOR_reg_22_inst : FD1 port map( D => n6673, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_22_port, QN => n_1422);
   KEY_EXPAN0_reg_63_22_inst : FD1 port map( D => n6061, CP => CLK_I, Q => 
                           n_1423, QN => n1291);
   KEY_EXPAN0_reg_62_22_inst : FD1 port map( D => n6060, CP => CLK_I, Q => 
                           n_1424, QN => n220);
   KEY_EXPAN0_reg_61_22_inst : FD1 port map( D => n6059, CP => CLK_I, Q => 
                           n_1425, QN => n1290);
   KEY_EXPAN0_reg_60_22_inst : FD1 port map( D => n6058, CP => CLK_I, Q => 
                           n_1426, QN => n219);
   KEY_EXPAN0_reg_59_22_inst : FD1 port map( D => n6057, CP => CLK_I, Q => 
                           n_1427, QN => n1289);
   KEY_EXPAN0_reg_58_22_inst : FD1 port map( D => n6056, CP => CLK_I, Q => 
                           n_1428, QN => n218);
   KEY_EXPAN0_reg_57_22_inst : FD1 port map( D => n6055, CP => CLK_I, Q => 
                           n_1429, QN => n1288);
   KEY_EXPAN0_reg_56_22_inst : FD1 port map( D => n6054, CP => CLK_I, Q => 
                           n_1430, QN => n217);
   KEY_EXPAN0_reg_55_22_inst : FD1 port map( D => n6053, CP => CLK_I, Q => 
                           n_1431, QN => n1295);
   KEY_EXPAN0_reg_54_22_inst : FD1 port map( D => n6052, CP => CLK_I, Q => 
                           n_1432, QN => n224);
   KEY_EXPAN0_reg_53_22_inst : FD1 port map( D => n6051, CP => CLK_I, Q => 
                           n_1433, QN => n1294);
   KEY_EXPAN0_reg_52_22_inst : FD1 port map( D => n6050, CP => CLK_I, Q => 
                           n_1434, QN => n223);
   KEY_EXPAN0_reg_51_22_inst : FD1 port map( D => n6049, CP => CLK_I, Q => 
                           n_1435, QN => n1293);
   KEY_EXPAN0_reg_50_22_inst : FD1 port map( D => n6048, CP => CLK_I, Q => 
                           n_1436, QN => n222);
   KEY_EXPAN0_reg_49_22_inst : FD1 port map( D => n6047, CP => CLK_I, Q => 
                           n_1437, QN => n1292);
   KEY_EXPAN0_reg_48_22_inst : FD1 port map( D => n6046, CP => CLK_I, Q => 
                           n_1438, QN => n221);
   KEY_EXPAN0_reg_47_22_inst : FD1 port map( D => n6045, CP => CLK_I, Q => 
                           n_1439, QN => n1299);
   KEY_EXPAN0_reg_46_22_inst : FD1 port map( D => n6044, CP => CLK_I, Q => 
                           n_1440, QN => n228);
   KEY_EXPAN0_reg_45_22_inst : FD1 port map( D => n6043, CP => CLK_I, Q => 
                           n_1441, QN => n1298);
   KEY_EXPAN0_reg_44_22_inst : FD1 port map( D => n6042, CP => CLK_I, Q => 
                           n_1442, QN => n227);
   KEY_EXPAN0_reg_43_22_inst : FD1 port map( D => n6041, CP => CLK_I, Q => 
                           n_1443, QN => n1297);
   KEY_EXPAN0_reg_42_22_inst : FD1 port map( D => n6040, CP => CLK_I, Q => 
                           n_1444, QN => n226);
   KEY_EXPAN0_reg_41_22_inst : FD1 port map( D => n6039, CP => CLK_I, Q => 
                           n_1445, QN => n1296);
   KEY_EXPAN0_reg_40_22_inst : FD1 port map( D => n6038, CP => CLK_I, Q => 
                           n_1446, QN => n225);
   KEY_EXPAN0_reg_39_22_inst : FD1 port map( D => n6037, CP => CLK_I, Q => 
                           n_1447, QN => n1303);
   KEY_EXPAN0_reg_38_22_inst : FD1 port map( D => n6036, CP => CLK_I, Q => 
                           n_1448, QN => n232);
   KEY_EXPAN0_reg_37_22_inst : FD1 port map( D => n6035, CP => CLK_I, Q => 
                           n_1449, QN => n1302);
   KEY_EXPAN0_reg_36_22_inst : FD1 port map( D => n6034, CP => CLK_I, Q => 
                           n_1450, QN => n231);
   KEY_EXPAN0_reg_35_22_inst : FD1 port map( D => n6033, CP => CLK_I, Q => 
                           n_1451, QN => n1301);
   KEY_EXPAN0_reg_34_22_inst : FD1 port map( D => n6032, CP => CLK_I, Q => 
                           n_1452, QN => n230);
   KEY_EXPAN0_reg_33_22_inst : FD1 port map( D => n6031, CP => CLK_I, Q => 
                           n_1453, QN => n1300);
   KEY_EXPAN0_reg_32_22_inst : FD1 port map( D => n6030, CP => CLK_I, Q => 
                           n_1454, QN => n229);
   KEY_EXPAN0_reg_31_22_inst : FD1 port map( D => n6029, CP => CLK_I, Q => 
                           n_1455, QN => n1275);
   KEY_EXPAN0_reg_30_22_inst : FD1 port map( D => n6028, CP => CLK_I, Q => 
                           n_1456, QN => n204);
   KEY_EXPAN0_reg_29_22_inst : FD1 port map( D => n6027, CP => CLK_I, Q => 
                           n_1457, QN => n1274);
   KEY_EXPAN0_reg_28_22_inst : FD1 port map( D => n6026, CP => CLK_I, Q => 
                           n_1458, QN => n203);
   KEY_EXPAN0_reg_27_22_inst : FD1 port map( D => n6025, CP => CLK_I, Q => 
                           n_1459, QN => n1273);
   KEY_EXPAN0_reg_26_22_inst : FD1 port map( D => n6024, CP => CLK_I, Q => 
                           n_1460, QN => n202);
   KEY_EXPAN0_reg_25_22_inst : FD1 port map( D => n6023, CP => CLK_I, Q => 
                           n_1461, QN => n1272);
   KEY_EXPAN0_reg_24_22_inst : FD1 port map( D => n6022, CP => CLK_I, Q => 
                           n_1462, QN => n201);
   KEY_EXPAN0_reg_23_22_inst : FD1 port map( D => n6021, CP => CLK_I, Q => 
                           n_1463, QN => n1279);
   KEY_EXPAN0_reg_22_22_inst : FD1 port map( D => n6020, CP => CLK_I, Q => 
                           n_1464, QN => n208);
   KEY_EXPAN0_reg_21_22_inst : FD1 port map( D => n6019, CP => CLK_I, Q => 
                           n_1465, QN => n1278);
   KEY_EXPAN0_reg_20_22_inst : FD1 port map( D => n6018, CP => CLK_I, Q => 
                           n_1466, QN => n207);
   KEY_EXPAN0_reg_19_22_inst : FD1 port map( D => n6017, CP => CLK_I, Q => 
                           n_1467, QN => n1277);
   KEY_EXPAN0_reg_18_22_inst : FD1 port map( D => n6016, CP => CLK_I, Q => 
                           n_1468, QN => n206);
   KEY_EXPAN0_reg_17_22_inst : FD1 port map( D => n6015, CP => CLK_I, Q => 
                           n_1469, QN => n1276);
   KEY_EXPAN0_reg_16_22_inst : FD1 port map( D => n6014, CP => CLK_I, Q => 
                           n_1470, QN => n205);
   KEY_EXPAN0_reg_15_22_inst : FD1 port map( D => n6013, CP => CLK_I, Q => 
                           n_1471, QN => n1283);
   KEY_EXPAN0_reg_14_22_inst : FD1 port map( D => n6012, CP => CLK_I, Q => 
                           n_1472, QN => n212);
   KEY_EXPAN0_reg_13_22_inst : FD1 port map( D => n6011, CP => CLK_I, Q => 
                           n_1473, QN => n1282);
   KEY_EXPAN0_reg_12_22_inst : FD1 port map( D => n6010, CP => CLK_I, Q => 
                           n_1474, QN => n211);
   KEY_EXPAN0_reg_11_22_inst : FD1 port map( D => n6009, CP => CLK_I, Q => 
                           n_1475, QN => n1281);
   KEY_EXPAN0_reg_10_22_inst : FD1 port map( D => n6008, CP => CLK_I, Q => 
                           n_1476, QN => n210);
   KEY_EXPAN0_reg_9_22_inst : FD1 port map( D => n6007, CP => CLK_I, Q => 
                           n_1477, QN => n1280);
   KEY_EXPAN0_reg_8_22_inst : FD1 port map( D => n6006, CP => CLK_I, Q => 
                           n_1478, QN => n209);
   KEY_EXPAN0_reg_7_22_inst : FD1 port map( D => n6005, CP => CLK_I, Q => 
                           n_1479, QN => n1287);
   KEY_EXPAN0_reg_6_22_inst : FD1 port map( D => n6004, CP => CLK_I, Q => 
                           n_1480, QN => n216);
   KEY_EXPAN0_reg_5_22_inst : FD1 port map( D => n6003, CP => CLK_I, Q => 
                           n_1481, QN => n1286);
   KEY_EXPAN0_reg_4_22_inst : FD1 port map( D => n6002, CP => CLK_I, Q => 
                           n_1482, QN => n215);
   KEY_EXPAN0_reg_3_22_inst : FD1 port map( D => n6001, CP => CLK_I, Q => 
                           n_1483, QN => n1285);
   KEY_EXPAN0_reg_2_22_inst : FD1 port map( D => n6000, CP => CLK_I, Q => 
                           n_1484, QN => n214);
   KEY_EXPAN0_reg_1_22_inst : FD1 port map( D => n5999, CP => CLK_I, Q => 
                           n_1485, QN => n1284);
   KEY_EXPAN0_reg_0_22_inst : FD1 port map( D => n5998, CP => CLK_I, Q => 
                           n_1486, QN => n213);
   v_KEY_COL_OUT0_reg_22_inst : FD1 port map( D => n4574, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_22_port, QN => n1060);
   v_TEMP_VECTOR_reg_14_inst : FD1 port map( D => n6681, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_14_port, QN => n_1487);
   KEY_EXPAN0_reg_63_14_inst : FD1 port map( D => n5549, CP => CLK_I, Q => 
                           n_1488, QN => n1323);
   KEY_EXPAN0_reg_62_14_inst : FD1 port map( D => n5548, CP => CLK_I, Q => 
                           n_1489, QN => n252);
   KEY_EXPAN0_reg_61_14_inst : FD1 port map( D => n5547, CP => CLK_I, Q => 
                           n_1490, QN => n1322);
   KEY_EXPAN0_reg_60_14_inst : FD1 port map( D => n5546, CP => CLK_I, Q => 
                           n_1491, QN => n251);
   KEY_EXPAN0_reg_59_14_inst : FD1 port map( D => n5545, CP => CLK_I, Q => 
                           n_1492, QN => n1321);
   KEY_EXPAN0_reg_58_14_inst : FD1 port map( D => n5544, CP => CLK_I, Q => 
                           n_1493, QN => n250);
   KEY_EXPAN0_reg_57_14_inst : FD1 port map( D => n5543, CP => CLK_I, Q => 
                           n_1494, QN => n1320);
   KEY_EXPAN0_reg_56_14_inst : FD1 port map( D => n5542, CP => CLK_I, Q => 
                           n_1495, QN => n249);
   KEY_EXPAN0_reg_55_14_inst : FD1 port map( D => n5541, CP => CLK_I, Q => 
                           n_1496, QN => n1327);
   KEY_EXPAN0_reg_54_14_inst : FD1 port map( D => n5540, CP => CLK_I, Q => 
                           n_1497, QN => n256);
   KEY_EXPAN0_reg_53_14_inst : FD1 port map( D => n5539, CP => CLK_I, Q => 
                           n_1498, QN => n1326);
   KEY_EXPAN0_reg_52_14_inst : FD1 port map( D => n5538, CP => CLK_I, Q => 
                           n_1499, QN => n255);
   KEY_EXPAN0_reg_51_14_inst : FD1 port map( D => n5537, CP => CLK_I, Q => 
                           n_1500, QN => n1325);
   KEY_EXPAN0_reg_50_14_inst : FD1 port map( D => n5536, CP => CLK_I, Q => 
                           n_1501, QN => n254);
   KEY_EXPAN0_reg_49_14_inst : FD1 port map( D => n5535, CP => CLK_I, Q => 
                           n_1502, QN => n1324);
   KEY_EXPAN0_reg_48_14_inst : FD1 port map( D => n5534, CP => CLK_I, Q => 
                           n_1503, QN => n253);
   KEY_EXPAN0_reg_47_14_inst : FD1 port map( D => n5533, CP => CLK_I, Q => 
                           n_1504, QN => n1331);
   KEY_EXPAN0_reg_46_14_inst : FD1 port map( D => n5532, CP => CLK_I, Q => 
                           n_1505, QN => n260);
   KEY_EXPAN0_reg_45_14_inst : FD1 port map( D => n5531, CP => CLK_I, Q => 
                           n_1506, QN => n1330);
   KEY_EXPAN0_reg_44_14_inst : FD1 port map( D => n5530, CP => CLK_I, Q => 
                           n_1507, QN => n259);
   KEY_EXPAN0_reg_43_14_inst : FD1 port map( D => n5529, CP => CLK_I, Q => 
                           n_1508, QN => n1329);
   KEY_EXPAN0_reg_42_14_inst : FD1 port map( D => n5528, CP => CLK_I, Q => 
                           n_1509, QN => n258);
   KEY_EXPAN0_reg_41_14_inst : FD1 port map( D => n5527, CP => CLK_I, Q => 
                           n_1510, QN => n1328);
   KEY_EXPAN0_reg_40_14_inst : FD1 port map( D => n5526, CP => CLK_I, Q => 
                           n_1511, QN => n257);
   KEY_EXPAN0_reg_39_14_inst : FD1 port map( D => n5525, CP => CLK_I, Q => 
                           n_1512, QN => n1335);
   KEY_EXPAN0_reg_38_14_inst : FD1 port map( D => n5524, CP => CLK_I, Q => 
                           n_1513, QN => n264);
   KEY_EXPAN0_reg_37_14_inst : FD1 port map( D => n5523, CP => CLK_I, Q => 
                           n_1514, QN => n1334);
   KEY_EXPAN0_reg_36_14_inst : FD1 port map( D => n5522, CP => CLK_I, Q => 
                           n_1515, QN => n263);
   KEY_EXPAN0_reg_35_14_inst : FD1 port map( D => n5521, CP => CLK_I, Q => 
                           n_1516, QN => n1333);
   KEY_EXPAN0_reg_34_14_inst : FD1 port map( D => n5520, CP => CLK_I, Q => 
                           n_1517, QN => n262);
   KEY_EXPAN0_reg_33_14_inst : FD1 port map( D => n5519, CP => CLK_I, Q => 
                           n_1518, QN => n1332);
   KEY_EXPAN0_reg_32_14_inst : FD1 port map( D => n5518, CP => CLK_I, Q => 
                           n_1519, QN => n261);
   KEY_EXPAN0_reg_31_14_inst : FD1 port map( D => n5517, CP => CLK_I, Q => 
                           n_1520, QN => n1307);
   KEY_EXPAN0_reg_30_14_inst : FD1 port map( D => n5516, CP => CLK_I, Q => 
                           n_1521, QN => n236);
   KEY_EXPAN0_reg_29_14_inst : FD1 port map( D => n5515, CP => CLK_I, Q => 
                           n_1522, QN => n1306);
   KEY_EXPAN0_reg_28_14_inst : FD1 port map( D => n5514, CP => CLK_I, Q => 
                           n_1523, QN => n235);
   KEY_EXPAN0_reg_27_14_inst : FD1 port map( D => n5513, CP => CLK_I, Q => 
                           n_1524, QN => n1305);
   KEY_EXPAN0_reg_26_14_inst : FD1 port map( D => n5512, CP => CLK_I, Q => 
                           n_1525, QN => n234);
   KEY_EXPAN0_reg_25_14_inst : FD1 port map( D => n5511, CP => CLK_I, Q => 
                           n_1526, QN => n1304);
   KEY_EXPAN0_reg_24_14_inst : FD1 port map( D => n5510, CP => CLK_I, Q => 
                           n_1527, QN => n233);
   KEY_EXPAN0_reg_23_14_inst : FD1 port map( D => n5509, CP => CLK_I, Q => 
                           n_1528, QN => n1311);
   KEY_EXPAN0_reg_22_14_inst : FD1 port map( D => n5508, CP => CLK_I, Q => 
                           n_1529, QN => n240);
   KEY_EXPAN0_reg_21_14_inst : FD1 port map( D => n5507, CP => CLK_I, Q => 
                           n_1530, QN => n1310);
   KEY_EXPAN0_reg_20_14_inst : FD1 port map( D => n5506, CP => CLK_I, Q => 
                           n_1531, QN => n239);
   KEY_EXPAN0_reg_19_14_inst : FD1 port map( D => n5505, CP => CLK_I, Q => 
                           n_1532, QN => n1309);
   KEY_EXPAN0_reg_18_14_inst : FD1 port map( D => n5504, CP => CLK_I, Q => 
                           n_1533, QN => n238);
   KEY_EXPAN0_reg_17_14_inst : FD1 port map( D => n5503, CP => CLK_I, Q => 
                           n_1534, QN => n1308);
   KEY_EXPAN0_reg_16_14_inst : FD1 port map( D => n5502, CP => CLK_I, Q => 
                           n_1535, QN => n237);
   KEY_EXPAN0_reg_15_14_inst : FD1 port map( D => n5501, CP => CLK_I, Q => 
                           n_1536, QN => n1315);
   KEY_EXPAN0_reg_14_14_inst : FD1 port map( D => n5500, CP => CLK_I, Q => 
                           n_1537, QN => n244);
   KEY_EXPAN0_reg_13_14_inst : FD1 port map( D => n5499, CP => CLK_I, Q => 
                           n_1538, QN => n1314);
   KEY_EXPAN0_reg_12_14_inst : FD1 port map( D => n5498, CP => CLK_I, Q => 
                           n_1539, QN => n243);
   KEY_EXPAN0_reg_11_14_inst : FD1 port map( D => n5497, CP => CLK_I, Q => 
                           n_1540, QN => n1313);
   KEY_EXPAN0_reg_10_14_inst : FD1 port map( D => n5496, CP => CLK_I, Q => 
                           n_1541, QN => n242);
   KEY_EXPAN0_reg_9_14_inst : FD1 port map( D => n5495, CP => CLK_I, Q => 
                           n_1542, QN => n1312);
   KEY_EXPAN0_reg_8_14_inst : FD1 port map( D => n5494, CP => CLK_I, Q => 
                           n_1543, QN => n241);
   KEY_EXPAN0_reg_7_14_inst : FD1 port map( D => n5493, CP => CLK_I, Q => 
                           n_1544, QN => n1319);
   KEY_EXPAN0_reg_6_14_inst : FD1 port map( D => n5492, CP => CLK_I, Q => 
                           n_1545, QN => n248);
   KEY_EXPAN0_reg_5_14_inst : FD1 port map( D => n5491, CP => CLK_I, Q => 
                           n_1546, QN => n1318);
   KEY_EXPAN0_reg_4_14_inst : FD1 port map( D => n5490, CP => CLK_I, Q => 
                           n_1547, QN => n247);
   KEY_EXPAN0_reg_3_14_inst : FD1 port map( D => n5489, CP => CLK_I, Q => 
                           n_1548, QN => n1317);
   KEY_EXPAN0_reg_2_14_inst : FD1 port map( D => n5488, CP => CLK_I, Q => 
                           n_1549, QN => n246);
   KEY_EXPAN0_reg_1_14_inst : FD1 port map( D => n5487, CP => CLK_I, Q => 
                           n_1550, QN => n1316);
   KEY_EXPAN0_reg_0_14_inst : FD1 port map( D => n5486, CP => CLK_I, Q => 
                           n_1551, QN => n245);
   v_KEY_COL_OUT0_reg_14_inst : FD1 port map( D => n4573, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_14_port, QN => n1069);
   v_TEMP_VECTOR_reg_5_inst : FD1 port map( D => n6690, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_5_port, QN => n_1552);
   KEY_EXPAN0_reg_63_5_inst : FD1 port map( D => n4973, CP => CLK_I, Q => 
                           n_1553, QN => n1355);
   KEY_EXPAN0_reg_62_5_inst : FD1 port map( D => n4972, CP => CLK_I, Q => 
                           n_1554, QN => n284);
   KEY_EXPAN0_reg_61_5_inst : FD1 port map( D => n4971, CP => CLK_I, Q => 
                           n_1555, QN => n1354);
   KEY_EXPAN0_reg_60_5_inst : FD1 port map( D => n4970, CP => CLK_I, Q => 
                           n_1556, QN => n283);
   KEY_EXPAN0_reg_59_5_inst : FD1 port map( D => n4969, CP => CLK_I, Q => 
                           n_1557, QN => n1353);
   KEY_EXPAN0_reg_58_5_inst : FD1 port map( D => n4968, CP => CLK_I, Q => 
                           n_1558, QN => n282);
   KEY_EXPAN0_reg_57_5_inst : FD1 port map( D => n4967, CP => CLK_I, Q => 
                           n_1559, QN => n1352);
   KEY_EXPAN0_reg_56_5_inst : FD1 port map( D => n4966, CP => CLK_I, Q => 
                           n_1560, QN => n281);
   KEY_EXPAN0_reg_55_5_inst : FD1 port map( D => n4965, CP => CLK_I, Q => 
                           n_1561, QN => n1359);
   KEY_EXPAN0_reg_54_5_inst : FD1 port map( D => n4964, CP => CLK_I, Q => 
                           n_1562, QN => n288);
   KEY_EXPAN0_reg_53_5_inst : FD1 port map( D => n4963, CP => CLK_I, Q => 
                           n_1563, QN => n1358);
   KEY_EXPAN0_reg_52_5_inst : FD1 port map( D => n4962, CP => CLK_I, Q => 
                           n_1564, QN => n287);
   KEY_EXPAN0_reg_51_5_inst : FD1 port map( D => n4961, CP => CLK_I, Q => 
                           n_1565, QN => n1357);
   KEY_EXPAN0_reg_50_5_inst : FD1 port map( D => n4960, CP => CLK_I, Q => 
                           n_1566, QN => n286);
   KEY_EXPAN0_reg_49_5_inst : FD1 port map( D => n4959, CP => CLK_I, Q => 
                           n_1567, QN => n1356);
   KEY_EXPAN0_reg_48_5_inst : FD1 port map( D => n4958, CP => CLK_I, Q => 
                           n_1568, QN => n285);
   KEY_EXPAN0_reg_47_5_inst : FD1 port map( D => n4957, CP => CLK_I, Q => 
                           n_1569, QN => n1363);
   KEY_EXPAN0_reg_46_5_inst : FD1 port map( D => n4956, CP => CLK_I, Q => 
                           n_1570, QN => n292);
   KEY_EXPAN0_reg_45_5_inst : FD1 port map( D => n4955, CP => CLK_I, Q => 
                           n_1571, QN => n1362);
   KEY_EXPAN0_reg_44_5_inst : FD1 port map( D => n4954, CP => CLK_I, Q => 
                           n_1572, QN => n291);
   KEY_EXPAN0_reg_43_5_inst : FD1 port map( D => n4953, CP => CLK_I, Q => 
                           n_1573, QN => n1361);
   KEY_EXPAN0_reg_42_5_inst : FD1 port map( D => n4952, CP => CLK_I, Q => 
                           n_1574, QN => n290);
   KEY_EXPAN0_reg_41_5_inst : FD1 port map( D => n4951, CP => CLK_I, Q => 
                           n_1575, QN => n1360);
   KEY_EXPAN0_reg_40_5_inst : FD1 port map( D => n4950, CP => CLK_I, Q => 
                           n_1576, QN => n289);
   KEY_EXPAN0_reg_39_5_inst : FD1 port map( D => n4949, CP => CLK_I, Q => 
                           n_1577, QN => n1367);
   KEY_EXPAN0_reg_38_5_inst : FD1 port map( D => n4948, CP => CLK_I, Q => 
                           n_1578, QN => n296);
   KEY_EXPAN0_reg_37_5_inst : FD1 port map( D => n4947, CP => CLK_I, Q => 
                           n_1579, QN => n1366);
   KEY_EXPAN0_reg_36_5_inst : FD1 port map( D => n4946, CP => CLK_I, Q => 
                           n_1580, QN => n295);
   KEY_EXPAN0_reg_35_5_inst : FD1 port map( D => n4945, CP => CLK_I, Q => 
                           n_1581, QN => n1365);
   KEY_EXPAN0_reg_34_5_inst : FD1 port map( D => n4944, CP => CLK_I, Q => 
                           n_1582, QN => n294);
   KEY_EXPAN0_reg_33_5_inst : FD1 port map( D => n4943, CP => CLK_I, Q => 
                           n_1583, QN => n1364);
   KEY_EXPAN0_reg_32_5_inst : FD1 port map( D => n4942, CP => CLK_I, Q => 
                           n_1584, QN => n293);
   KEY_EXPAN0_reg_31_5_inst : FD1 port map( D => n4941, CP => CLK_I, Q => 
                           n_1585, QN => n1339);
   KEY_EXPAN0_reg_30_5_inst : FD1 port map( D => n4940, CP => CLK_I, Q => 
                           n_1586, QN => n268);
   KEY_EXPAN0_reg_29_5_inst : FD1 port map( D => n4939, CP => CLK_I, Q => 
                           n_1587, QN => n1338);
   KEY_EXPAN0_reg_28_5_inst : FD1 port map( D => n4938, CP => CLK_I, Q => 
                           n_1588, QN => n267);
   KEY_EXPAN0_reg_27_5_inst : FD1 port map( D => n4937, CP => CLK_I, Q => 
                           n_1589, QN => n1337);
   KEY_EXPAN0_reg_26_5_inst : FD1 port map( D => n4936, CP => CLK_I, Q => 
                           n_1590, QN => n266);
   KEY_EXPAN0_reg_25_5_inst : FD1 port map( D => n4935, CP => CLK_I, Q => 
                           n_1591, QN => n1336);
   KEY_EXPAN0_reg_24_5_inst : FD1 port map( D => n4934, CP => CLK_I, Q => 
                           n_1592, QN => n265);
   KEY_EXPAN0_reg_23_5_inst : FD1 port map( D => n4933, CP => CLK_I, Q => 
                           n_1593, QN => n1343);
   KEY_EXPAN0_reg_22_5_inst : FD1 port map( D => n4932, CP => CLK_I, Q => 
                           n_1594, QN => n272);
   KEY_EXPAN0_reg_21_5_inst : FD1 port map( D => n4931, CP => CLK_I, Q => 
                           n_1595, QN => n1342);
   KEY_EXPAN0_reg_20_5_inst : FD1 port map( D => n4930, CP => CLK_I, Q => 
                           n_1596, QN => n271);
   KEY_EXPAN0_reg_19_5_inst : FD1 port map( D => n4929, CP => CLK_I, Q => 
                           n_1597, QN => n1341);
   KEY_EXPAN0_reg_18_5_inst : FD1 port map( D => n4928, CP => CLK_I, Q => 
                           n_1598, QN => n270);
   KEY_EXPAN0_reg_17_5_inst : FD1 port map( D => n4927, CP => CLK_I, Q => 
                           n_1599, QN => n1340);
   KEY_EXPAN0_reg_16_5_inst : FD1 port map( D => n4926, CP => CLK_I, Q => 
                           n_1600, QN => n269);
   KEY_EXPAN0_reg_15_5_inst : FD1 port map( D => n4925, CP => CLK_I, Q => 
                           n_1601, QN => n1347);
   KEY_EXPAN0_reg_14_5_inst : FD1 port map( D => n4924, CP => CLK_I, Q => 
                           n_1602, QN => n276);
   KEY_EXPAN0_reg_13_5_inst : FD1 port map( D => n4923, CP => CLK_I, Q => 
                           n_1603, QN => n1346);
   KEY_EXPAN0_reg_12_5_inst : FD1 port map( D => n4922, CP => CLK_I, Q => 
                           n_1604, QN => n275);
   KEY_EXPAN0_reg_11_5_inst : FD1 port map( D => n4921, CP => CLK_I, Q => 
                           n_1605, QN => n1345);
   KEY_EXPAN0_reg_10_5_inst : FD1 port map( D => n4920, CP => CLK_I, Q => 
                           n_1606, QN => n274);
   KEY_EXPAN0_reg_9_5_inst : FD1 port map( D => n4919, CP => CLK_I, Q => n_1607
                           , QN => n1344);
   KEY_EXPAN0_reg_8_5_inst : FD1 port map( D => n4918, CP => CLK_I, Q => n_1608
                           , QN => n273);
   KEY_EXPAN0_reg_7_5_inst : FD1 port map( D => n4917, CP => CLK_I, Q => n_1609
                           , QN => n1351);
   KEY_EXPAN0_reg_6_5_inst : FD1 port map( D => n4916, CP => CLK_I, Q => n_1610
                           , QN => n280);
   KEY_EXPAN0_reg_5_5_inst : FD1 port map( D => n4915, CP => CLK_I, Q => n_1611
                           , QN => n1350);
   KEY_EXPAN0_reg_4_5_inst : FD1 port map( D => n4914, CP => CLK_I, Q => n_1612
                           , QN => n279);
   KEY_EXPAN0_reg_3_5_inst : FD1 port map( D => n4913, CP => CLK_I, Q => n_1613
                           , QN => n1349);
   KEY_EXPAN0_reg_2_5_inst : FD1 port map( D => n4912, CP => CLK_I, Q => n_1614
                           , QN => n278);
   KEY_EXPAN0_reg_1_5_inst : FD1 port map( D => n4911, CP => CLK_I, Q => n_1615
                           , QN => n1348);
   KEY_EXPAN0_reg_0_5_inst : FD1 port map( D => n4910, CP => CLK_I, Q => n_1616
                           , QN => n277);
   v_KEY_COL_OUT0_reg_5_inst : FD1 port map( D => n4572, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_5_port, QN => n1047);
   v_TEMP_VECTOR_reg_29_inst : FD1 port map( D => n6666, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_29_port, QN => n_1617);
   KEY_EXPAN0_reg_63_29_inst : FD1 port map( D => n6509, CP => CLK_I, Q => 
                           n_1618, QN => n1387);
   KEY_EXPAN0_reg_62_29_inst : FD1 port map( D => n6508, CP => CLK_I, Q => 
                           n_1619, QN => n316);
   KEY_EXPAN0_reg_61_29_inst : FD1 port map( D => n6507, CP => CLK_I, Q => 
                           n_1620, QN => n1386);
   KEY_EXPAN0_reg_60_29_inst : FD1 port map( D => n6506, CP => CLK_I, Q => 
                           n_1621, QN => n315);
   KEY_EXPAN0_reg_59_29_inst : FD1 port map( D => n6505, CP => CLK_I, Q => 
                           n_1622, QN => n1385);
   KEY_EXPAN0_reg_58_29_inst : FD1 port map( D => n6504, CP => CLK_I, Q => 
                           n_1623, QN => n314);
   KEY_EXPAN0_reg_57_29_inst : FD1 port map( D => n6503, CP => CLK_I, Q => 
                           n_1624, QN => n1384);
   KEY_EXPAN0_reg_56_29_inst : FD1 port map( D => n6502, CP => CLK_I, Q => 
                           n_1625, QN => n313);
   KEY_EXPAN0_reg_55_29_inst : FD1 port map( D => n6501, CP => CLK_I, Q => 
                           n_1626, QN => n1391);
   KEY_EXPAN0_reg_54_29_inst : FD1 port map( D => n6500, CP => CLK_I, Q => 
                           n_1627, QN => n320);
   KEY_EXPAN0_reg_53_29_inst : FD1 port map( D => n6499, CP => CLK_I, Q => 
                           n_1628, QN => n1390);
   KEY_EXPAN0_reg_52_29_inst : FD1 port map( D => n6498, CP => CLK_I, Q => 
                           n_1629, QN => n319);
   KEY_EXPAN0_reg_51_29_inst : FD1 port map( D => n6497, CP => CLK_I, Q => 
                           n_1630, QN => n1389);
   KEY_EXPAN0_reg_50_29_inst : FD1 port map( D => n6496, CP => CLK_I, Q => 
                           n_1631, QN => n318);
   KEY_EXPAN0_reg_49_29_inst : FD1 port map( D => n6495, CP => CLK_I, Q => 
                           n_1632, QN => n1388);
   KEY_EXPAN0_reg_48_29_inst : FD1 port map( D => n6494, CP => CLK_I, Q => 
                           n_1633, QN => n317);
   KEY_EXPAN0_reg_47_29_inst : FD1 port map( D => n6493, CP => CLK_I, Q => 
                           n_1634, QN => n1395);
   KEY_EXPAN0_reg_46_29_inst : FD1 port map( D => n6492, CP => CLK_I, Q => 
                           n_1635, QN => n324);
   KEY_EXPAN0_reg_45_29_inst : FD1 port map( D => n6491, CP => CLK_I, Q => 
                           n_1636, QN => n1394);
   KEY_EXPAN0_reg_44_29_inst : FD1 port map( D => n6490, CP => CLK_I, Q => 
                           n_1637, QN => n323);
   KEY_EXPAN0_reg_43_29_inst : FD1 port map( D => n6489, CP => CLK_I, Q => 
                           n_1638, QN => n1393);
   KEY_EXPAN0_reg_42_29_inst : FD1 port map( D => n6488, CP => CLK_I, Q => 
                           n_1639, QN => n322);
   KEY_EXPAN0_reg_41_29_inst : FD1 port map( D => n6487, CP => CLK_I, Q => 
                           n_1640, QN => n1392);
   KEY_EXPAN0_reg_40_29_inst : FD1 port map( D => n6486, CP => CLK_I, Q => 
                           n_1641, QN => n321);
   KEY_EXPAN0_reg_39_29_inst : FD1 port map( D => n6485, CP => CLK_I, Q => 
                           n_1642, QN => n1399);
   KEY_EXPAN0_reg_38_29_inst : FD1 port map( D => n6484, CP => CLK_I, Q => 
                           n_1643, QN => n328);
   KEY_EXPAN0_reg_37_29_inst : FD1 port map( D => n6483, CP => CLK_I, Q => 
                           n_1644, QN => n1398);
   KEY_EXPAN0_reg_36_29_inst : FD1 port map( D => n6482, CP => CLK_I, Q => 
                           n_1645, QN => n327);
   KEY_EXPAN0_reg_35_29_inst : FD1 port map( D => n6481, CP => CLK_I, Q => 
                           n_1646, QN => n1397);
   KEY_EXPAN0_reg_34_29_inst : FD1 port map( D => n6480, CP => CLK_I, Q => 
                           n_1647, QN => n326);
   KEY_EXPAN0_reg_33_29_inst : FD1 port map( D => n6479, CP => CLK_I, Q => 
                           n_1648, QN => n1396);
   KEY_EXPAN0_reg_32_29_inst : FD1 port map( D => n6478, CP => CLK_I, Q => 
                           n_1649, QN => n325);
   KEY_EXPAN0_reg_31_29_inst : FD1 port map( D => n6477, CP => CLK_I, Q => 
                           n_1650, QN => n1371);
   KEY_EXPAN0_reg_30_29_inst : FD1 port map( D => n6476, CP => CLK_I, Q => 
                           n_1651, QN => n300);
   KEY_EXPAN0_reg_29_29_inst : FD1 port map( D => n6475, CP => CLK_I, Q => 
                           n_1652, QN => n1370);
   KEY_EXPAN0_reg_28_29_inst : FD1 port map( D => n6474, CP => CLK_I, Q => 
                           n_1653, QN => n299);
   KEY_EXPAN0_reg_27_29_inst : FD1 port map( D => n6473, CP => CLK_I, Q => 
                           n_1654, QN => n1369);
   KEY_EXPAN0_reg_26_29_inst : FD1 port map( D => n6472, CP => CLK_I, Q => 
                           n_1655, QN => n298);
   KEY_EXPAN0_reg_25_29_inst : FD1 port map( D => n6471, CP => CLK_I, Q => 
                           n_1656, QN => n1368);
   KEY_EXPAN0_reg_24_29_inst : FD1 port map( D => n6470, CP => CLK_I, Q => 
                           n_1657, QN => n297);
   KEY_EXPAN0_reg_23_29_inst : FD1 port map( D => n6469, CP => CLK_I, Q => 
                           n_1658, QN => n1375);
   KEY_EXPAN0_reg_22_29_inst : FD1 port map( D => n6468, CP => CLK_I, Q => 
                           n_1659, QN => n304);
   KEY_EXPAN0_reg_21_29_inst : FD1 port map( D => n6467, CP => CLK_I, Q => 
                           n_1660, QN => n1374);
   KEY_EXPAN0_reg_20_29_inst : FD1 port map( D => n6466, CP => CLK_I, Q => 
                           n_1661, QN => n303);
   KEY_EXPAN0_reg_19_29_inst : FD1 port map( D => n6465, CP => CLK_I, Q => 
                           n_1662, QN => n1373);
   KEY_EXPAN0_reg_18_29_inst : FD1 port map( D => n6464, CP => CLK_I, Q => 
                           n_1663, QN => n302);
   KEY_EXPAN0_reg_17_29_inst : FD1 port map( D => n6463, CP => CLK_I, Q => 
                           n_1664, QN => n1372);
   KEY_EXPAN0_reg_16_29_inst : FD1 port map( D => n6462, CP => CLK_I, Q => 
                           n_1665, QN => n301);
   KEY_EXPAN0_reg_15_29_inst : FD1 port map( D => n6461, CP => CLK_I, Q => 
                           n_1666, QN => n1379);
   KEY_EXPAN0_reg_14_29_inst : FD1 port map( D => n6460, CP => CLK_I, Q => 
                           n_1667, QN => n308);
   KEY_EXPAN0_reg_13_29_inst : FD1 port map( D => n6459, CP => CLK_I, Q => 
                           n_1668, QN => n1378);
   KEY_EXPAN0_reg_12_29_inst : FD1 port map( D => n6458, CP => CLK_I, Q => 
                           n_1669, QN => n307);
   KEY_EXPAN0_reg_11_29_inst : FD1 port map( D => n6457, CP => CLK_I, Q => 
                           n_1670, QN => n1377);
   KEY_EXPAN0_reg_10_29_inst : FD1 port map( D => n6456, CP => CLK_I, Q => 
                           n_1671, QN => n306);
   KEY_EXPAN0_reg_9_29_inst : FD1 port map( D => n6455, CP => CLK_I, Q => 
                           n_1672, QN => n1376);
   KEY_EXPAN0_reg_8_29_inst : FD1 port map( D => n6454, CP => CLK_I, Q => 
                           n_1673, QN => n305);
   KEY_EXPAN0_reg_7_29_inst : FD1 port map( D => n6453, CP => CLK_I, Q => 
                           n_1674, QN => n1383);
   KEY_EXPAN0_reg_6_29_inst : FD1 port map( D => n6452, CP => CLK_I, Q => 
                           n_1675, QN => n312);
   KEY_EXPAN0_reg_5_29_inst : FD1 port map( D => n6451, CP => CLK_I, Q => 
                           n_1676, QN => n1382);
   KEY_EXPAN0_reg_4_29_inst : FD1 port map( D => n6450, CP => CLK_I, Q => 
                           n_1677, QN => n311);
   KEY_EXPAN0_reg_3_29_inst : FD1 port map( D => n6449, CP => CLK_I, Q => 
                           n_1678, QN => n1381);
   KEY_EXPAN0_reg_2_29_inst : FD1 port map( D => n6448, CP => CLK_I, Q => 
                           n_1679, QN => n310);
   KEY_EXPAN0_reg_1_29_inst : FD1 port map( D => n6447, CP => CLK_I, Q => 
                           n_1680, QN => n1380);
   KEY_EXPAN0_reg_0_29_inst : FD1 port map( D => n6446, CP => CLK_I, Q => 
                           n_1681, QN => n309);
   v_KEY_COL_OUT0_reg_29_inst : FD1 port map( D => n4571, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_29_port, QN => n1053);
   v_TEMP_VECTOR_reg_21_inst : FD1 port map( D => n6674, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_21_port, QN => n_1682);
   KEY_EXPAN0_reg_63_21_inst : FD1 port map( D => n5997, CP => CLK_I, Q => 
                           n_1683, QN => n1419);
   KEY_EXPAN0_reg_62_21_inst : FD1 port map( D => n5996, CP => CLK_I, Q => 
                           n_1684, QN => n348);
   KEY_EXPAN0_reg_61_21_inst : FD1 port map( D => n5995, CP => CLK_I, Q => 
                           n_1685, QN => n1418);
   KEY_EXPAN0_reg_60_21_inst : FD1 port map( D => n5994, CP => CLK_I, Q => 
                           n_1686, QN => n347);
   KEY_EXPAN0_reg_59_21_inst : FD1 port map( D => n5993, CP => CLK_I, Q => 
                           n_1687, QN => n1417);
   KEY_EXPAN0_reg_58_21_inst : FD1 port map( D => n5992, CP => CLK_I, Q => 
                           n_1688, QN => n346);
   KEY_EXPAN0_reg_57_21_inst : FD1 port map( D => n5991, CP => CLK_I, Q => 
                           n_1689, QN => n1416);
   KEY_EXPAN0_reg_56_21_inst : FD1 port map( D => n5990, CP => CLK_I, Q => 
                           n_1690, QN => n345);
   KEY_EXPAN0_reg_55_21_inst : FD1 port map( D => n5989, CP => CLK_I, Q => 
                           n_1691, QN => n1423);
   KEY_EXPAN0_reg_54_21_inst : FD1 port map( D => n5988, CP => CLK_I, Q => 
                           n_1692, QN => n352);
   KEY_EXPAN0_reg_53_21_inst : FD1 port map( D => n5987, CP => CLK_I, Q => 
                           n_1693, QN => n1422);
   KEY_EXPAN0_reg_52_21_inst : FD1 port map( D => n5986, CP => CLK_I, Q => 
                           n_1694, QN => n351);
   KEY_EXPAN0_reg_51_21_inst : FD1 port map( D => n5985, CP => CLK_I, Q => 
                           n_1695, QN => n1421);
   KEY_EXPAN0_reg_50_21_inst : FD1 port map( D => n5984, CP => CLK_I, Q => 
                           n_1696, QN => n350);
   KEY_EXPAN0_reg_49_21_inst : FD1 port map( D => n5983, CP => CLK_I, Q => 
                           n_1697, QN => n1420);
   KEY_EXPAN0_reg_48_21_inst : FD1 port map( D => n5982, CP => CLK_I, Q => 
                           n_1698, QN => n349);
   KEY_EXPAN0_reg_47_21_inst : FD1 port map( D => n5981, CP => CLK_I, Q => 
                           n_1699, QN => n1427);
   KEY_EXPAN0_reg_46_21_inst : FD1 port map( D => n5980, CP => CLK_I, Q => 
                           n_1700, QN => n356);
   KEY_EXPAN0_reg_45_21_inst : FD1 port map( D => n5979, CP => CLK_I, Q => 
                           n_1701, QN => n1426);
   KEY_EXPAN0_reg_44_21_inst : FD1 port map( D => n5978, CP => CLK_I, Q => 
                           n_1702, QN => n355);
   KEY_EXPAN0_reg_43_21_inst : FD1 port map( D => n5977, CP => CLK_I, Q => 
                           n_1703, QN => n1425);
   KEY_EXPAN0_reg_42_21_inst : FD1 port map( D => n5976, CP => CLK_I, Q => 
                           n_1704, QN => n354);
   KEY_EXPAN0_reg_41_21_inst : FD1 port map( D => n5975, CP => CLK_I, Q => 
                           n_1705, QN => n1424);
   KEY_EXPAN0_reg_40_21_inst : FD1 port map( D => n5974, CP => CLK_I, Q => 
                           n_1706, QN => n353);
   KEY_EXPAN0_reg_39_21_inst : FD1 port map( D => n5973, CP => CLK_I, Q => 
                           n_1707, QN => n1431);
   KEY_EXPAN0_reg_38_21_inst : FD1 port map( D => n5972, CP => CLK_I, Q => 
                           n_1708, QN => n360);
   KEY_EXPAN0_reg_37_21_inst : FD1 port map( D => n5971, CP => CLK_I, Q => 
                           n_1709, QN => n1430);
   KEY_EXPAN0_reg_36_21_inst : FD1 port map( D => n5970, CP => CLK_I, Q => 
                           n_1710, QN => n359);
   KEY_EXPAN0_reg_35_21_inst : FD1 port map( D => n5969, CP => CLK_I, Q => 
                           n_1711, QN => n1429);
   KEY_EXPAN0_reg_34_21_inst : FD1 port map( D => n5968, CP => CLK_I, Q => 
                           n_1712, QN => n358);
   KEY_EXPAN0_reg_33_21_inst : FD1 port map( D => n5967, CP => CLK_I, Q => 
                           n_1713, QN => n1428);
   KEY_EXPAN0_reg_32_21_inst : FD1 port map( D => n5966, CP => CLK_I, Q => 
                           n_1714, QN => n357);
   KEY_EXPAN0_reg_31_21_inst : FD1 port map( D => n5965, CP => CLK_I, Q => 
                           n_1715, QN => n1403);
   KEY_EXPAN0_reg_30_21_inst : FD1 port map( D => n5964, CP => CLK_I, Q => 
                           n_1716, QN => n332);
   KEY_EXPAN0_reg_29_21_inst : FD1 port map( D => n5963, CP => CLK_I, Q => 
                           n_1717, QN => n1402);
   KEY_EXPAN0_reg_28_21_inst : FD1 port map( D => n5962, CP => CLK_I, Q => 
                           n_1718, QN => n331);
   KEY_EXPAN0_reg_27_21_inst : FD1 port map( D => n5961, CP => CLK_I, Q => 
                           n_1719, QN => n1401);
   KEY_EXPAN0_reg_26_21_inst : FD1 port map( D => n5960, CP => CLK_I, Q => 
                           n_1720, QN => n330);
   KEY_EXPAN0_reg_25_21_inst : FD1 port map( D => n5959, CP => CLK_I, Q => 
                           n_1721, QN => n1400);
   KEY_EXPAN0_reg_24_21_inst : FD1 port map( D => n5958, CP => CLK_I, Q => 
                           n_1722, QN => n329);
   KEY_EXPAN0_reg_23_21_inst : FD1 port map( D => n5957, CP => CLK_I, Q => 
                           n_1723, QN => n1407);
   KEY_EXPAN0_reg_22_21_inst : FD1 port map( D => n5956, CP => CLK_I, Q => 
                           n_1724, QN => n336);
   KEY_EXPAN0_reg_21_21_inst : FD1 port map( D => n5955, CP => CLK_I, Q => 
                           n_1725, QN => n1406);
   KEY_EXPAN0_reg_20_21_inst : FD1 port map( D => n5954, CP => CLK_I, Q => 
                           n_1726, QN => n335);
   KEY_EXPAN0_reg_19_21_inst : FD1 port map( D => n5953, CP => CLK_I, Q => 
                           n_1727, QN => n1405);
   KEY_EXPAN0_reg_18_21_inst : FD1 port map( D => n5952, CP => CLK_I, Q => 
                           n_1728, QN => n334);
   KEY_EXPAN0_reg_17_21_inst : FD1 port map( D => n5951, CP => CLK_I, Q => 
                           n_1729, QN => n1404);
   KEY_EXPAN0_reg_16_21_inst : FD1 port map( D => n5950, CP => CLK_I, Q => 
                           n_1730, QN => n333);
   KEY_EXPAN0_reg_15_21_inst : FD1 port map( D => n5949, CP => CLK_I, Q => 
                           n_1731, QN => n1411);
   KEY_EXPAN0_reg_14_21_inst : FD1 port map( D => n5948, CP => CLK_I, Q => 
                           n_1732, QN => n340);
   KEY_EXPAN0_reg_13_21_inst : FD1 port map( D => n5947, CP => CLK_I, Q => 
                           n_1733, QN => n1410);
   KEY_EXPAN0_reg_12_21_inst : FD1 port map( D => n5946, CP => CLK_I, Q => 
                           n_1734, QN => n339);
   KEY_EXPAN0_reg_11_21_inst : FD1 port map( D => n5945, CP => CLK_I, Q => 
                           n_1735, QN => n1409);
   KEY_EXPAN0_reg_10_21_inst : FD1 port map( D => n5944, CP => CLK_I, Q => 
                           n_1736, QN => n338);
   KEY_EXPAN0_reg_9_21_inst : FD1 port map( D => n5943, CP => CLK_I, Q => 
                           n_1737, QN => n1408);
   KEY_EXPAN0_reg_8_21_inst : FD1 port map( D => n5942, CP => CLK_I, Q => 
                           n_1738, QN => n337);
   KEY_EXPAN0_reg_7_21_inst : FD1 port map( D => n5941, CP => CLK_I, Q => 
                           n_1739, QN => n1415);
   KEY_EXPAN0_reg_6_21_inst : FD1 port map( D => n5940, CP => CLK_I, Q => 
                           n_1740, QN => n344);
   KEY_EXPAN0_reg_5_21_inst : FD1 port map( D => n5939, CP => CLK_I, Q => 
                           n_1741, QN => n1414);
   KEY_EXPAN0_reg_4_21_inst : FD1 port map( D => n5938, CP => CLK_I, Q => 
                           n_1742, QN => n343);
   KEY_EXPAN0_reg_3_21_inst : FD1 port map( D => n5937, CP => CLK_I, Q => 
                           n_1743, QN => n1413);
   KEY_EXPAN0_reg_2_21_inst : FD1 port map( D => n5936, CP => CLK_I, Q => 
                           n_1744, QN => n342);
   KEY_EXPAN0_reg_1_21_inst : FD1 port map( D => n5935, CP => CLK_I, Q => 
                           n_1745, QN => n1412);
   KEY_EXPAN0_reg_0_21_inst : FD1 port map( D => n5934, CP => CLK_I, Q => 
                           n_1746, QN => n341);
   v_KEY_COL_OUT0_reg_21_inst : FD1 port map( D => n4570, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_21_port, QN => n1061);
   v_TEMP_VECTOR_reg_13_inst : FD1 port map( D => n6682, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_13_port, QN => n_1747);
   KEY_EXPAN0_reg_63_13_inst : FD1 port map( D => n5485, CP => CLK_I, Q => 
                           n_1748, QN => n1451);
   KEY_EXPAN0_reg_62_13_inst : FD1 port map( D => n5484, CP => CLK_I, Q => 
                           n_1749, QN => n380);
   KEY_EXPAN0_reg_61_13_inst : FD1 port map( D => n5483, CP => CLK_I, Q => 
                           n_1750, QN => n1450);
   KEY_EXPAN0_reg_60_13_inst : FD1 port map( D => n5482, CP => CLK_I, Q => 
                           n_1751, QN => n379);
   KEY_EXPAN0_reg_59_13_inst : FD1 port map( D => n5481, CP => CLK_I, Q => 
                           n_1752, QN => n1449);
   KEY_EXPAN0_reg_58_13_inst : FD1 port map( D => n5480, CP => CLK_I, Q => 
                           n_1753, QN => n378);
   KEY_EXPAN0_reg_57_13_inst : FD1 port map( D => n5479, CP => CLK_I, Q => 
                           n_1754, QN => n1448);
   KEY_EXPAN0_reg_56_13_inst : FD1 port map( D => n5478, CP => CLK_I, Q => 
                           n_1755, QN => n377);
   KEY_EXPAN0_reg_55_13_inst : FD1 port map( D => n5477, CP => CLK_I, Q => 
                           n_1756, QN => n1455);
   KEY_EXPAN0_reg_54_13_inst : FD1 port map( D => n5476, CP => CLK_I, Q => 
                           n_1757, QN => n384);
   KEY_EXPAN0_reg_53_13_inst : FD1 port map( D => n5475, CP => CLK_I, Q => 
                           n_1758, QN => n1454);
   KEY_EXPAN0_reg_52_13_inst : FD1 port map( D => n5474, CP => CLK_I, Q => 
                           n_1759, QN => n383);
   KEY_EXPAN0_reg_51_13_inst : FD1 port map( D => n5473, CP => CLK_I, Q => 
                           n_1760, QN => n1453);
   KEY_EXPAN0_reg_50_13_inst : FD1 port map( D => n5472, CP => CLK_I, Q => 
                           n_1761, QN => n382);
   KEY_EXPAN0_reg_49_13_inst : FD1 port map( D => n5471, CP => CLK_I, Q => 
                           n_1762, QN => n1452);
   KEY_EXPAN0_reg_48_13_inst : FD1 port map( D => n5470, CP => CLK_I, Q => 
                           n_1763, QN => n381);
   KEY_EXPAN0_reg_47_13_inst : FD1 port map( D => n5469, CP => CLK_I, Q => 
                           n_1764, QN => n1459);
   KEY_EXPAN0_reg_46_13_inst : FD1 port map( D => n5468, CP => CLK_I, Q => 
                           n_1765, QN => n388);
   KEY_EXPAN0_reg_45_13_inst : FD1 port map( D => n5467, CP => CLK_I, Q => 
                           n_1766, QN => n1458);
   KEY_EXPAN0_reg_44_13_inst : FD1 port map( D => n5466, CP => CLK_I, Q => 
                           n_1767, QN => n387);
   KEY_EXPAN0_reg_43_13_inst : FD1 port map( D => n5465, CP => CLK_I, Q => 
                           n_1768, QN => n1457);
   KEY_EXPAN0_reg_42_13_inst : FD1 port map( D => n5464, CP => CLK_I, Q => 
                           n_1769, QN => n386);
   KEY_EXPAN0_reg_41_13_inst : FD1 port map( D => n5463, CP => CLK_I, Q => 
                           n_1770, QN => n1456);
   KEY_EXPAN0_reg_40_13_inst : FD1 port map( D => n5462, CP => CLK_I, Q => 
                           n_1771, QN => n385);
   KEY_EXPAN0_reg_39_13_inst : FD1 port map( D => n5461, CP => CLK_I, Q => 
                           n_1772, QN => n1463);
   KEY_EXPAN0_reg_38_13_inst : FD1 port map( D => n5460, CP => CLK_I, Q => 
                           n_1773, QN => n392);
   KEY_EXPAN0_reg_37_13_inst : FD1 port map( D => n5459, CP => CLK_I, Q => 
                           n_1774, QN => n1462);
   KEY_EXPAN0_reg_36_13_inst : FD1 port map( D => n5458, CP => CLK_I, Q => 
                           n_1775, QN => n391);
   KEY_EXPAN0_reg_35_13_inst : FD1 port map( D => n5457, CP => CLK_I, Q => 
                           n_1776, QN => n1461);
   KEY_EXPAN0_reg_34_13_inst : FD1 port map( D => n5456, CP => CLK_I, Q => 
                           n_1777, QN => n390);
   KEY_EXPAN0_reg_33_13_inst : FD1 port map( D => n5455, CP => CLK_I, Q => 
                           n_1778, QN => n1460);
   KEY_EXPAN0_reg_32_13_inst : FD1 port map( D => n5454, CP => CLK_I, Q => 
                           n_1779, QN => n389);
   KEY_EXPAN0_reg_31_13_inst : FD1 port map( D => n5453, CP => CLK_I, Q => 
                           n_1780, QN => n1435);
   KEY_EXPAN0_reg_30_13_inst : FD1 port map( D => n5452, CP => CLK_I, Q => 
                           n_1781, QN => n364);
   KEY_EXPAN0_reg_29_13_inst : FD1 port map( D => n5451, CP => CLK_I, Q => 
                           n_1782, QN => n1434);
   KEY_EXPAN0_reg_28_13_inst : FD1 port map( D => n5450, CP => CLK_I, Q => 
                           n_1783, QN => n363);
   KEY_EXPAN0_reg_27_13_inst : FD1 port map( D => n5449, CP => CLK_I, Q => 
                           n_1784, QN => n1433);
   KEY_EXPAN0_reg_26_13_inst : FD1 port map( D => n5448, CP => CLK_I, Q => 
                           n_1785, QN => n362);
   KEY_EXPAN0_reg_25_13_inst : FD1 port map( D => n5447, CP => CLK_I, Q => 
                           n_1786, QN => n1432);
   KEY_EXPAN0_reg_24_13_inst : FD1 port map( D => n5446, CP => CLK_I, Q => 
                           n_1787, QN => n361);
   KEY_EXPAN0_reg_23_13_inst : FD1 port map( D => n5445, CP => CLK_I, Q => 
                           n_1788, QN => n1439);
   KEY_EXPAN0_reg_22_13_inst : FD1 port map( D => n5444, CP => CLK_I, Q => 
                           n_1789, QN => n368);
   KEY_EXPAN0_reg_21_13_inst : FD1 port map( D => n5443, CP => CLK_I, Q => 
                           n_1790, QN => n1438);
   KEY_EXPAN0_reg_20_13_inst : FD1 port map( D => n5442, CP => CLK_I, Q => 
                           n_1791, QN => n367);
   KEY_EXPAN0_reg_19_13_inst : FD1 port map( D => n5441, CP => CLK_I, Q => 
                           n_1792, QN => n1437);
   KEY_EXPAN0_reg_18_13_inst : FD1 port map( D => n5440, CP => CLK_I, Q => 
                           n_1793, QN => n366);
   KEY_EXPAN0_reg_17_13_inst : FD1 port map( D => n5439, CP => CLK_I, Q => 
                           n_1794, QN => n1436);
   KEY_EXPAN0_reg_16_13_inst : FD1 port map( D => n5438, CP => CLK_I, Q => 
                           n_1795, QN => n365);
   KEY_EXPAN0_reg_15_13_inst : FD1 port map( D => n5437, CP => CLK_I, Q => 
                           n_1796, QN => n1443);
   KEY_EXPAN0_reg_14_13_inst : FD1 port map( D => n5436, CP => CLK_I, Q => 
                           n_1797, QN => n372);
   KEY_EXPAN0_reg_13_13_inst : FD1 port map( D => n5435, CP => CLK_I, Q => 
                           n_1798, QN => n1442);
   KEY_EXPAN0_reg_12_13_inst : FD1 port map( D => n5434, CP => CLK_I, Q => 
                           n_1799, QN => n371);
   KEY_EXPAN0_reg_11_13_inst : FD1 port map( D => n5433, CP => CLK_I, Q => 
                           n_1800, QN => n1441);
   KEY_EXPAN0_reg_10_13_inst : FD1 port map( D => n5432, CP => CLK_I, Q => 
                           n_1801, QN => n370);
   KEY_EXPAN0_reg_9_13_inst : FD1 port map( D => n5431, CP => CLK_I, Q => 
                           n_1802, QN => n1440);
   KEY_EXPAN0_reg_8_13_inst : FD1 port map( D => n5430, CP => CLK_I, Q => 
                           n_1803, QN => n369);
   KEY_EXPAN0_reg_7_13_inst : FD1 port map( D => n5429, CP => CLK_I, Q => 
                           n_1804, QN => n1447);
   KEY_EXPAN0_reg_6_13_inst : FD1 port map( D => n5428, CP => CLK_I, Q => 
                           n_1805, QN => n376);
   KEY_EXPAN0_reg_5_13_inst : FD1 port map( D => n5427, CP => CLK_I, Q => 
                           n_1806, QN => n1446);
   KEY_EXPAN0_reg_4_13_inst : FD1 port map( D => n5426, CP => CLK_I, Q => 
                           n_1807, QN => n375);
   KEY_EXPAN0_reg_3_13_inst : FD1 port map( D => n5425, CP => CLK_I, Q => 
                           n_1808, QN => n1445);
   KEY_EXPAN0_reg_2_13_inst : FD1 port map( D => n5424, CP => CLK_I, Q => 
                           n_1809, QN => n374);
   KEY_EXPAN0_reg_1_13_inst : FD1 port map( D => n5423, CP => CLK_I, Q => 
                           n_1810, QN => n1444);
   KEY_EXPAN0_reg_0_13_inst : FD1 port map( D => n5422, CP => CLK_I, Q => 
                           n_1811, QN => n373);
   v_KEY_COL_OUT0_reg_13_inst : FD1 port map( D => n4569, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_13_port, QN => n1070);
   v_TEMP_VECTOR_reg_4_inst : FD1 port map( D => n6691, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_4_port, QN => n_1812);
   KEY_EXPAN0_reg_63_4_inst : FD1 port map( D => n4909, CP => CLK_I, Q => 
                           n_1813, QN => n1483);
   KEY_EXPAN0_reg_62_4_inst : FD1 port map( D => n4908, CP => CLK_I, Q => 
                           n_1814, QN => n412);
   KEY_EXPAN0_reg_61_4_inst : FD1 port map( D => n4907, CP => CLK_I, Q => 
                           n_1815, QN => n1482);
   KEY_EXPAN0_reg_60_4_inst : FD1 port map( D => n4906, CP => CLK_I, Q => 
                           n_1816, QN => n411);
   KEY_EXPAN0_reg_59_4_inst : FD1 port map( D => n4905, CP => CLK_I, Q => 
                           n_1817, QN => n1481);
   KEY_EXPAN0_reg_58_4_inst : FD1 port map( D => n4904, CP => CLK_I, Q => 
                           n_1818, QN => n410);
   KEY_EXPAN0_reg_57_4_inst : FD1 port map( D => n4903, CP => CLK_I, Q => 
                           n_1819, QN => n1480);
   KEY_EXPAN0_reg_56_4_inst : FD1 port map( D => n4902, CP => CLK_I, Q => 
                           n_1820, QN => n409);
   KEY_EXPAN0_reg_55_4_inst : FD1 port map( D => n4901, CP => CLK_I, Q => 
                           n_1821, QN => n1487);
   KEY_EXPAN0_reg_54_4_inst : FD1 port map( D => n4900, CP => CLK_I, Q => 
                           n_1822, QN => n416);
   KEY_EXPAN0_reg_53_4_inst : FD1 port map( D => n4899, CP => CLK_I, Q => 
                           n_1823, QN => n1486);
   KEY_EXPAN0_reg_52_4_inst : FD1 port map( D => n4898, CP => CLK_I, Q => 
                           n_1824, QN => n415);
   KEY_EXPAN0_reg_51_4_inst : FD1 port map( D => n4897, CP => CLK_I, Q => 
                           n_1825, QN => n1485);
   KEY_EXPAN0_reg_50_4_inst : FD1 port map( D => n4896, CP => CLK_I, Q => 
                           n_1826, QN => n414);
   KEY_EXPAN0_reg_49_4_inst : FD1 port map( D => n4895, CP => CLK_I, Q => 
                           n_1827, QN => n1484);
   KEY_EXPAN0_reg_48_4_inst : FD1 port map( D => n4894, CP => CLK_I, Q => 
                           n_1828, QN => n413);
   KEY_EXPAN0_reg_47_4_inst : FD1 port map( D => n4893, CP => CLK_I, Q => 
                           n_1829, QN => n1491);
   KEY_EXPAN0_reg_46_4_inst : FD1 port map( D => n4892, CP => CLK_I, Q => 
                           n_1830, QN => n420);
   KEY_EXPAN0_reg_45_4_inst : FD1 port map( D => n4891, CP => CLK_I, Q => 
                           n_1831, QN => n1490);
   KEY_EXPAN0_reg_44_4_inst : FD1 port map( D => n4890, CP => CLK_I, Q => 
                           n_1832, QN => n419);
   KEY_EXPAN0_reg_43_4_inst : FD1 port map( D => n4889, CP => CLK_I, Q => 
                           n_1833, QN => n1489);
   KEY_EXPAN0_reg_42_4_inst : FD1 port map( D => n4888, CP => CLK_I, Q => 
                           n_1834, QN => n418);
   KEY_EXPAN0_reg_41_4_inst : FD1 port map( D => n4887, CP => CLK_I, Q => 
                           n_1835, QN => n1488);
   KEY_EXPAN0_reg_40_4_inst : FD1 port map( D => n4886, CP => CLK_I, Q => 
                           n_1836, QN => n417);
   KEY_EXPAN0_reg_39_4_inst : FD1 port map( D => n4885, CP => CLK_I, Q => 
                           n_1837, QN => n1495);
   KEY_EXPAN0_reg_38_4_inst : FD1 port map( D => n4884, CP => CLK_I, Q => 
                           n_1838, QN => n424);
   KEY_EXPAN0_reg_37_4_inst : FD1 port map( D => n4883, CP => CLK_I, Q => 
                           n_1839, QN => n1494);
   KEY_EXPAN0_reg_36_4_inst : FD1 port map( D => n4882, CP => CLK_I, Q => 
                           n_1840, QN => n423);
   KEY_EXPAN0_reg_35_4_inst : FD1 port map( D => n4881, CP => CLK_I, Q => 
                           n_1841, QN => n1493);
   KEY_EXPAN0_reg_34_4_inst : FD1 port map( D => n4880, CP => CLK_I, Q => 
                           n_1842, QN => n422);
   KEY_EXPAN0_reg_33_4_inst : FD1 port map( D => n4879, CP => CLK_I, Q => 
                           n_1843, QN => n1492);
   KEY_EXPAN0_reg_32_4_inst : FD1 port map( D => n4878, CP => CLK_I, Q => 
                           n_1844, QN => n421);
   KEY_EXPAN0_reg_31_4_inst : FD1 port map( D => n4877, CP => CLK_I, Q => 
                           n_1845, QN => n1467);
   KEY_EXPAN0_reg_30_4_inst : FD1 port map( D => n4876, CP => CLK_I, Q => 
                           n_1846, QN => n396);
   KEY_EXPAN0_reg_29_4_inst : FD1 port map( D => n4875, CP => CLK_I, Q => 
                           n_1847, QN => n1466);
   KEY_EXPAN0_reg_28_4_inst : FD1 port map( D => n4874, CP => CLK_I, Q => 
                           n_1848, QN => n395);
   KEY_EXPAN0_reg_27_4_inst : FD1 port map( D => n4873, CP => CLK_I, Q => 
                           n_1849, QN => n1465);
   KEY_EXPAN0_reg_26_4_inst : FD1 port map( D => n4872, CP => CLK_I, Q => 
                           n_1850, QN => n394);
   KEY_EXPAN0_reg_25_4_inst : FD1 port map( D => n4871, CP => CLK_I, Q => 
                           n_1851, QN => n1464);
   KEY_EXPAN0_reg_24_4_inst : FD1 port map( D => n4870, CP => CLK_I, Q => 
                           n_1852, QN => n393);
   KEY_EXPAN0_reg_23_4_inst : FD1 port map( D => n4869, CP => CLK_I, Q => 
                           n_1853, QN => n1471);
   KEY_EXPAN0_reg_22_4_inst : FD1 port map( D => n4868, CP => CLK_I, Q => 
                           n_1854, QN => n400);
   KEY_EXPAN0_reg_21_4_inst : FD1 port map( D => n4867, CP => CLK_I, Q => 
                           n_1855, QN => n1470);
   KEY_EXPAN0_reg_20_4_inst : FD1 port map( D => n4866, CP => CLK_I, Q => 
                           n_1856, QN => n399);
   KEY_EXPAN0_reg_19_4_inst : FD1 port map( D => n4865, CP => CLK_I, Q => 
                           n_1857, QN => n1469);
   KEY_EXPAN0_reg_18_4_inst : FD1 port map( D => n4864, CP => CLK_I, Q => 
                           n_1858, QN => n398);
   KEY_EXPAN0_reg_17_4_inst : FD1 port map( D => n4863, CP => CLK_I, Q => 
                           n_1859, QN => n1468);
   KEY_EXPAN0_reg_16_4_inst : FD1 port map( D => n4862, CP => CLK_I, Q => 
                           n_1860, QN => n397);
   KEY_EXPAN0_reg_15_4_inst : FD1 port map( D => n4861, CP => CLK_I, Q => 
                           n_1861, QN => n1475);
   KEY_EXPAN0_reg_14_4_inst : FD1 port map( D => n4860, CP => CLK_I, Q => 
                           n_1862, QN => n404);
   KEY_EXPAN0_reg_13_4_inst : FD1 port map( D => n4859, CP => CLK_I, Q => 
                           n_1863, QN => n1474);
   KEY_EXPAN0_reg_12_4_inst : FD1 port map( D => n4858, CP => CLK_I, Q => 
                           n_1864, QN => n403);
   KEY_EXPAN0_reg_11_4_inst : FD1 port map( D => n4857, CP => CLK_I, Q => 
                           n_1865, QN => n1473);
   KEY_EXPAN0_reg_10_4_inst : FD1 port map( D => n4856, CP => CLK_I, Q => 
                           n_1866, QN => n402);
   KEY_EXPAN0_reg_9_4_inst : FD1 port map( D => n4855, CP => CLK_I, Q => n_1867
                           , QN => n1472);
   KEY_EXPAN0_reg_8_4_inst : FD1 port map( D => n4854, CP => CLK_I, Q => n_1868
                           , QN => n401);
   KEY_EXPAN0_reg_7_4_inst : FD1 port map( D => n4853, CP => CLK_I, Q => n_1869
                           , QN => n1479);
   KEY_EXPAN0_reg_6_4_inst : FD1 port map( D => n4852, CP => CLK_I, Q => n_1870
                           , QN => n408);
   KEY_EXPAN0_reg_5_4_inst : FD1 port map( D => n4851, CP => CLK_I, Q => n_1871
                           , QN => n1478);
   KEY_EXPAN0_reg_4_4_inst : FD1 port map( D => n4850, CP => CLK_I, Q => n_1872
                           , QN => n407);
   KEY_EXPAN0_reg_3_4_inst : FD1 port map( D => n4849, CP => CLK_I, Q => n_1873
                           , QN => n1477);
   KEY_EXPAN0_reg_2_4_inst : FD1 port map( D => n4848, CP => CLK_I, Q => n_1874
                           , QN => n406);
   KEY_EXPAN0_reg_1_4_inst : FD1 port map( D => n4847, CP => CLK_I, Q => n_1875
                           , QN => n1476);
   KEY_EXPAN0_reg_0_4_inst : FD1 port map( D => n4846, CP => CLK_I, Q => n_1876
                           , QN => n405);
   v_KEY_COL_OUT0_reg_4_inst : FD1 port map( D => n4568, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_4_port, QN => n1048);
   v_TEMP_VECTOR_reg_28_inst : FD1 port map( D => n6667, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_28_port, QN => n_1877);
   KEY_EXPAN0_reg_63_28_inst : FD1 port map( D => n6445, CP => CLK_I, Q => 
                           n_1878, QN => n1515);
   KEY_EXPAN0_reg_62_28_inst : FD1 port map( D => n6444, CP => CLK_I, Q => 
                           n_1879, QN => n444);
   KEY_EXPAN0_reg_61_28_inst : FD1 port map( D => n6443, CP => CLK_I, Q => 
                           n_1880, QN => n1514);
   KEY_EXPAN0_reg_60_28_inst : FD1 port map( D => n6442, CP => CLK_I, Q => 
                           n_1881, QN => n443);
   KEY_EXPAN0_reg_59_28_inst : FD1 port map( D => n6441, CP => CLK_I, Q => 
                           n_1882, QN => n1513);
   KEY_EXPAN0_reg_58_28_inst : FD1 port map( D => n6440, CP => CLK_I, Q => 
                           n_1883, QN => n442);
   KEY_EXPAN0_reg_57_28_inst : FD1 port map( D => n6439, CP => CLK_I, Q => 
                           n_1884, QN => n1512);
   KEY_EXPAN0_reg_56_28_inst : FD1 port map( D => n6438, CP => CLK_I, Q => 
                           n_1885, QN => n441);
   KEY_EXPAN0_reg_55_28_inst : FD1 port map( D => n6437, CP => CLK_I, Q => 
                           n_1886, QN => n1519);
   KEY_EXPAN0_reg_54_28_inst : FD1 port map( D => n6436, CP => CLK_I, Q => 
                           n_1887, QN => n448);
   KEY_EXPAN0_reg_53_28_inst : FD1 port map( D => n6435, CP => CLK_I, Q => 
                           n_1888, QN => n1518);
   KEY_EXPAN0_reg_52_28_inst : FD1 port map( D => n6434, CP => CLK_I, Q => 
                           n_1889, QN => n447);
   KEY_EXPAN0_reg_51_28_inst : FD1 port map( D => n6433, CP => CLK_I, Q => 
                           n_1890, QN => n1517);
   KEY_EXPAN0_reg_50_28_inst : FD1 port map( D => n6432, CP => CLK_I, Q => 
                           n_1891, QN => n446);
   KEY_EXPAN0_reg_49_28_inst : FD1 port map( D => n6431, CP => CLK_I, Q => 
                           n_1892, QN => n1516);
   KEY_EXPAN0_reg_48_28_inst : FD1 port map( D => n6430, CP => CLK_I, Q => 
                           n_1893, QN => n445);
   KEY_EXPAN0_reg_47_28_inst : FD1 port map( D => n6429, CP => CLK_I, Q => 
                           n_1894, QN => n1523);
   KEY_EXPAN0_reg_46_28_inst : FD1 port map( D => n6428, CP => CLK_I, Q => 
                           n_1895, QN => n452);
   KEY_EXPAN0_reg_45_28_inst : FD1 port map( D => n6427, CP => CLK_I, Q => 
                           n_1896, QN => n1522);
   KEY_EXPAN0_reg_44_28_inst : FD1 port map( D => n6426, CP => CLK_I, Q => 
                           n_1897, QN => n451);
   KEY_EXPAN0_reg_43_28_inst : FD1 port map( D => n6425, CP => CLK_I, Q => 
                           n_1898, QN => n1521);
   KEY_EXPAN0_reg_42_28_inst : FD1 port map( D => n6424, CP => CLK_I, Q => 
                           n_1899, QN => n450);
   KEY_EXPAN0_reg_41_28_inst : FD1 port map( D => n6423, CP => CLK_I, Q => 
                           n_1900, QN => n1520);
   KEY_EXPAN0_reg_40_28_inst : FD1 port map( D => n6422, CP => CLK_I, Q => 
                           n_1901, QN => n449);
   KEY_EXPAN0_reg_39_28_inst : FD1 port map( D => n6421, CP => CLK_I, Q => 
                           n_1902, QN => n1527);
   KEY_EXPAN0_reg_38_28_inst : FD1 port map( D => n6420, CP => CLK_I, Q => 
                           n_1903, QN => n456);
   KEY_EXPAN0_reg_37_28_inst : FD1 port map( D => n6419, CP => CLK_I, Q => 
                           n_1904, QN => n1526);
   KEY_EXPAN0_reg_36_28_inst : FD1 port map( D => n6418, CP => CLK_I, Q => 
                           n_1905, QN => n455);
   KEY_EXPAN0_reg_35_28_inst : FD1 port map( D => n6417, CP => CLK_I, Q => 
                           n_1906, QN => n1525);
   KEY_EXPAN0_reg_34_28_inst : FD1 port map( D => n6416, CP => CLK_I, Q => 
                           n_1907, QN => n454);
   KEY_EXPAN0_reg_33_28_inst : FD1 port map( D => n6415, CP => CLK_I, Q => 
                           n_1908, QN => n1524);
   KEY_EXPAN0_reg_32_28_inst : FD1 port map( D => n6414, CP => CLK_I, Q => 
                           n_1909, QN => n453);
   KEY_EXPAN0_reg_31_28_inst : FD1 port map( D => n6413, CP => CLK_I, Q => 
                           n_1910, QN => n1499);
   KEY_EXPAN0_reg_30_28_inst : FD1 port map( D => n6412, CP => CLK_I, Q => 
                           n_1911, QN => n428);
   KEY_EXPAN0_reg_29_28_inst : FD1 port map( D => n6411, CP => CLK_I, Q => 
                           n_1912, QN => n1498);
   KEY_EXPAN0_reg_28_28_inst : FD1 port map( D => n6410, CP => CLK_I, Q => 
                           n_1913, QN => n427);
   KEY_EXPAN0_reg_27_28_inst : FD1 port map( D => n6409, CP => CLK_I, Q => 
                           n_1914, QN => n1497);
   KEY_EXPAN0_reg_26_28_inst : FD1 port map( D => n6408, CP => CLK_I, Q => 
                           n_1915, QN => n426);
   KEY_EXPAN0_reg_25_28_inst : FD1 port map( D => n6407, CP => CLK_I, Q => 
                           n_1916, QN => n1496);
   KEY_EXPAN0_reg_24_28_inst : FD1 port map( D => n6406, CP => CLK_I, Q => 
                           n_1917, QN => n425);
   KEY_EXPAN0_reg_23_28_inst : FD1 port map( D => n6405, CP => CLK_I, Q => 
                           n_1918, QN => n1503);
   KEY_EXPAN0_reg_22_28_inst : FD1 port map( D => n6404, CP => CLK_I, Q => 
                           n_1919, QN => n432);
   KEY_EXPAN0_reg_21_28_inst : FD1 port map( D => n6403, CP => CLK_I, Q => 
                           n_1920, QN => n1502);
   KEY_EXPAN0_reg_20_28_inst : FD1 port map( D => n6402, CP => CLK_I, Q => 
                           n_1921, QN => n431);
   KEY_EXPAN0_reg_19_28_inst : FD1 port map( D => n6401, CP => CLK_I, Q => 
                           n_1922, QN => n1501);
   KEY_EXPAN0_reg_18_28_inst : FD1 port map( D => n6400, CP => CLK_I, Q => 
                           n_1923, QN => n430);
   KEY_EXPAN0_reg_17_28_inst : FD1 port map( D => n6399, CP => CLK_I, Q => 
                           n_1924, QN => n1500);
   KEY_EXPAN0_reg_16_28_inst : FD1 port map( D => n6398, CP => CLK_I, Q => 
                           n_1925, QN => n429);
   KEY_EXPAN0_reg_15_28_inst : FD1 port map( D => n6397, CP => CLK_I, Q => 
                           n_1926, QN => n1507);
   KEY_EXPAN0_reg_14_28_inst : FD1 port map( D => n6396, CP => CLK_I, Q => 
                           n_1927, QN => n436);
   KEY_EXPAN0_reg_13_28_inst : FD1 port map( D => n6395, CP => CLK_I, Q => 
                           n_1928, QN => n1506);
   KEY_EXPAN0_reg_12_28_inst : FD1 port map( D => n6394, CP => CLK_I, Q => 
                           n_1929, QN => n435);
   KEY_EXPAN0_reg_11_28_inst : FD1 port map( D => n6393, CP => CLK_I, Q => 
                           n_1930, QN => n1505);
   KEY_EXPAN0_reg_10_28_inst : FD1 port map( D => n6392, CP => CLK_I, Q => 
                           n_1931, QN => n434);
   KEY_EXPAN0_reg_9_28_inst : FD1 port map( D => n6391, CP => CLK_I, Q => 
                           n_1932, QN => n1504);
   KEY_EXPAN0_reg_8_28_inst : FD1 port map( D => n6390, CP => CLK_I, Q => 
                           n_1933, QN => n433);
   KEY_EXPAN0_reg_7_28_inst : FD1 port map( D => n6389, CP => CLK_I, Q => 
                           n_1934, QN => n1511);
   KEY_EXPAN0_reg_6_28_inst : FD1 port map( D => n6388, CP => CLK_I, Q => 
                           n_1935, QN => n440);
   KEY_EXPAN0_reg_5_28_inst : FD1 port map( D => n6387, CP => CLK_I, Q => 
                           n_1936, QN => n1510);
   KEY_EXPAN0_reg_4_28_inst : FD1 port map( D => n6386, CP => CLK_I, Q => 
                           n_1937, QN => n439);
   KEY_EXPAN0_reg_3_28_inst : FD1 port map( D => n6385, CP => CLK_I, Q => 
                           n_1938, QN => n1509);
   KEY_EXPAN0_reg_2_28_inst : FD1 port map( D => n6384, CP => CLK_I, Q => 
                           n_1939, QN => n438);
   KEY_EXPAN0_reg_1_28_inst : FD1 port map( D => n6383, CP => CLK_I, Q => 
                           n_1940, QN => n1508);
   KEY_EXPAN0_reg_0_28_inst : FD1 port map( D => n6382, CP => CLK_I, Q => 
                           n_1941, QN => n437);
   v_KEY_COL_OUT0_reg_28_inst : FD1 port map( D => n4567, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_28_port, QN => n1054);
   v_TEMP_VECTOR_reg_20_inst : FD1 port map( D => n6675, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_20_port, QN => n_1942);
   KEY_EXPAN0_reg_63_20_inst : FD1 port map( D => n5933, CP => CLK_I, Q => 
                           n_1943, QN => n1547);
   KEY_EXPAN0_reg_62_20_inst : FD1 port map( D => n5932, CP => CLK_I, Q => 
                           n_1944, QN => n476);
   KEY_EXPAN0_reg_61_20_inst : FD1 port map( D => n5931, CP => CLK_I, Q => 
                           n_1945, QN => n1546);
   KEY_EXPAN0_reg_60_20_inst : FD1 port map( D => n5930, CP => CLK_I, Q => 
                           n_1946, QN => n475);
   KEY_EXPAN0_reg_59_20_inst : FD1 port map( D => n5929, CP => CLK_I, Q => 
                           n_1947, QN => n1545);
   KEY_EXPAN0_reg_58_20_inst : FD1 port map( D => n5928, CP => CLK_I, Q => 
                           n_1948, QN => n474);
   KEY_EXPAN0_reg_57_20_inst : FD1 port map( D => n5927, CP => CLK_I, Q => 
                           n_1949, QN => n1544);
   KEY_EXPAN0_reg_56_20_inst : FD1 port map( D => n5926, CP => CLK_I, Q => 
                           n_1950, QN => n473);
   KEY_EXPAN0_reg_55_20_inst : FD1 port map( D => n5925, CP => CLK_I, Q => 
                           n_1951, QN => n1551);
   KEY_EXPAN0_reg_54_20_inst : FD1 port map( D => n5924, CP => CLK_I, Q => 
                           n_1952, QN => n480);
   KEY_EXPAN0_reg_53_20_inst : FD1 port map( D => n5923, CP => CLK_I, Q => 
                           n_1953, QN => n1550);
   KEY_EXPAN0_reg_52_20_inst : FD1 port map( D => n5922, CP => CLK_I, Q => 
                           n_1954, QN => n479);
   KEY_EXPAN0_reg_51_20_inst : FD1 port map( D => n5921, CP => CLK_I, Q => 
                           n_1955, QN => n1549);
   KEY_EXPAN0_reg_50_20_inst : FD1 port map( D => n5920, CP => CLK_I, Q => 
                           n_1956, QN => n478);
   KEY_EXPAN0_reg_49_20_inst : FD1 port map( D => n5919, CP => CLK_I, Q => 
                           n_1957, QN => n1548);
   KEY_EXPAN0_reg_48_20_inst : FD1 port map( D => n5918, CP => CLK_I, Q => 
                           n_1958, QN => n477);
   KEY_EXPAN0_reg_47_20_inst : FD1 port map( D => n5917, CP => CLK_I, Q => 
                           n_1959, QN => n1555);
   KEY_EXPAN0_reg_46_20_inst : FD1 port map( D => n5916, CP => CLK_I, Q => 
                           n_1960, QN => n484);
   KEY_EXPAN0_reg_45_20_inst : FD1 port map( D => n5915, CP => CLK_I, Q => 
                           n_1961, QN => n1554);
   KEY_EXPAN0_reg_44_20_inst : FD1 port map( D => n5914, CP => CLK_I, Q => 
                           n_1962, QN => n483);
   KEY_EXPAN0_reg_43_20_inst : FD1 port map( D => n5913, CP => CLK_I, Q => 
                           n_1963, QN => n1553);
   KEY_EXPAN0_reg_42_20_inst : FD1 port map( D => n5912, CP => CLK_I, Q => 
                           n_1964, QN => n482);
   KEY_EXPAN0_reg_41_20_inst : FD1 port map( D => n5911, CP => CLK_I, Q => 
                           n_1965, QN => n1552);
   KEY_EXPAN0_reg_40_20_inst : FD1 port map( D => n5910, CP => CLK_I, Q => 
                           n_1966, QN => n481);
   KEY_EXPAN0_reg_39_20_inst : FD1 port map( D => n5909, CP => CLK_I, Q => 
                           n_1967, QN => n1559);
   KEY_EXPAN0_reg_38_20_inst : FD1 port map( D => n5908, CP => CLK_I, Q => 
                           n_1968, QN => n488);
   KEY_EXPAN0_reg_37_20_inst : FD1 port map( D => n5907, CP => CLK_I, Q => 
                           n_1969, QN => n1558);
   KEY_EXPAN0_reg_36_20_inst : FD1 port map( D => n5906, CP => CLK_I, Q => 
                           n_1970, QN => n487);
   KEY_EXPAN0_reg_35_20_inst : FD1 port map( D => n5905, CP => CLK_I, Q => 
                           n_1971, QN => n1557);
   KEY_EXPAN0_reg_34_20_inst : FD1 port map( D => n5904, CP => CLK_I, Q => 
                           n_1972, QN => n486);
   KEY_EXPAN0_reg_33_20_inst : FD1 port map( D => n5903, CP => CLK_I, Q => 
                           n_1973, QN => n1556);
   KEY_EXPAN0_reg_32_20_inst : FD1 port map( D => n5902, CP => CLK_I, Q => 
                           n_1974, QN => n485);
   KEY_EXPAN0_reg_31_20_inst : FD1 port map( D => n5901, CP => CLK_I, Q => 
                           n_1975, QN => n1531);
   KEY_EXPAN0_reg_30_20_inst : FD1 port map( D => n5900, CP => CLK_I, Q => 
                           n_1976, QN => n460);
   KEY_EXPAN0_reg_29_20_inst : FD1 port map( D => n5899, CP => CLK_I, Q => 
                           n_1977, QN => n1530);
   KEY_EXPAN0_reg_28_20_inst : FD1 port map( D => n5898, CP => CLK_I, Q => 
                           n_1978, QN => n459);
   KEY_EXPAN0_reg_27_20_inst : FD1 port map( D => n5897, CP => CLK_I, Q => 
                           n_1979, QN => n1529);
   KEY_EXPAN0_reg_26_20_inst : FD1 port map( D => n5896, CP => CLK_I, Q => 
                           n_1980, QN => n458);
   KEY_EXPAN0_reg_25_20_inst : FD1 port map( D => n5895, CP => CLK_I, Q => 
                           n_1981, QN => n1528);
   KEY_EXPAN0_reg_24_20_inst : FD1 port map( D => n5894, CP => CLK_I, Q => 
                           n_1982, QN => n457);
   KEY_EXPAN0_reg_23_20_inst : FD1 port map( D => n5893, CP => CLK_I, Q => 
                           n_1983, QN => n1535);
   KEY_EXPAN0_reg_22_20_inst : FD1 port map( D => n5892, CP => CLK_I, Q => 
                           n_1984, QN => n464);
   KEY_EXPAN0_reg_21_20_inst : FD1 port map( D => n5891, CP => CLK_I, Q => 
                           n_1985, QN => n1534);
   KEY_EXPAN0_reg_20_20_inst : FD1 port map( D => n5890, CP => CLK_I, Q => 
                           n_1986, QN => n463);
   KEY_EXPAN0_reg_19_20_inst : FD1 port map( D => n5889, CP => CLK_I, Q => 
                           n_1987, QN => n1533);
   KEY_EXPAN0_reg_18_20_inst : FD1 port map( D => n5888, CP => CLK_I, Q => 
                           n_1988, QN => n462);
   KEY_EXPAN0_reg_17_20_inst : FD1 port map( D => n5887, CP => CLK_I, Q => 
                           n_1989, QN => n1532);
   KEY_EXPAN0_reg_16_20_inst : FD1 port map( D => n5886, CP => CLK_I, Q => 
                           n_1990, QN => n461);
   KEY_EXPAN0_reg_15_20_inst : FD1 port map( D => n5885, CP => CLK_I, Q => 
                           n_1991, QN => n1539);
   KEY_EXPAN0_reg_14_20_inst : FD1 port map( D => n5884, CP => CLK_I, Q => 
                           n_1992, QN => n468);
   KEY_EXPAN0_reg_13_20_inst : FD1 port map( D => n5883, CP => CLK_I, Q => 
                           n_1993, QN => n1538);
   KEY_EXPAN0_reg_12_20_inst : FD1 port map( D => n5882, CP => CLK_I, Q => 
                           n_1994, QN => n467);
   KEY_EXPAN0_reg_11_20_inst : FD1 port map( D => n5881, CP => CLK_I, Q => 
                           n_1995, QN => n1537);
   KEY_EXPAN0_reg_10_20_inst : FD1 port map( D => n5880, CP => CLK_I, Q => 
                           n_1996, QN => n466);
   KEY_EXPAN0_reg_9_20_inst : FD1 port map( D => n5879, CP => CLK_I, Q => 
                           n_1997, QN => n1536);
   KEY_EXPAN0_reg_8_20_inst : FD1 port map( D => n5878, CP => CLK_I, Q => 
                           n_1998, QN => n465);
   KEY_EXPAN0_reg_7_20_inst : FD1 port map( D => n5877, CP => CLK_I, Q => 
                           n_1999, QN => n1543);
   KEY_EXPAN0_reg_6_20_inst : FD1 port map( D => n5876, CP => CLK_I, Q => 
                           n_2000, QN => n472);
   KEY_EXPAN0_reg_5_20_inst : FD1 port map( D => n5875, CP => CLK_I, Q => 
                           n_2001, QN => n1542);
   KEY_EXPAN0_reg_4_20_inst : FD1 port map( D => n5874, CP => CLK_I, Q => 
                           n_2002, QN => n471);
   KEY_EXPAN0_reg_3_20_inst : FD1 port map( D => n5873, CP => CLK_I, Q => 
                           n_2003, QN => n1541);
   KEY_EXPAN0_reg_2_20_inst : FD1 port map( D => n5872, CP => CLK_I, Q => 
                           n_2004, QN => n470);
   KEY_EXPAN0_reg_1_20_inst : FD1 port map( D => n5871, CP => CLK_I, Q => 
                           n_2005, QN => n1540);
   KEY_EXPAN0_reg_0_20_inst : FD1 port map( D => n5870, CP => CLK_I, Q => 
                           n_2006, QN => n469);
   v_KEY_COL_OUT0_reg_20_inst : FD1 port map( D => n4566, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_20_port, QN => n1062);
   v_TEMP_VECTOR_reg_12_inst : FD1 port map( D => n6683, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_12_port, QN => n_2007);
   KEY_EXPAN0_reg_63_12_inst : FD1 port map( D => n5421, CP => CLK_I, Q => 
                           n_2008, QN => n1579);
   KEY_EXPAN0_reg_62_12_inst : FD1 port map( D => n5420, CP => CLK_I, Q => 
                           n_2009, QN => n508);
   KEY_EXPAN0_reg_61_12_inst : FD1 port map( D => n5419, CP => CLK_I, Q => 
                           n_2010, QN => n1578);
   KEY_EXPAN0_reg_60_12_inst : FD1 port map( D => n5418, CP => CLK_I, Q => 
                           n_2011, QN => n507);
   KEY_EXPAN0_reg_59_12_inst : FD1 port map( D => n5417, CP => CLK_I, Q => 
                           n_2012, QN => n1577);
   KEY_EXPAN0_reg_58_12_inst : FD1 port map( D => n5416, CP => CLK_I, Q => 
                           n_2013, QN => n506);
   KEY_EXPAN0_reg_57_12_inst : FD1 port map( D => n5415, CP => CLK_I, Q => 
                           n_2014, QN => n1576);
   KEY_EXPAN0_reg_56_12_inst : FD1 port map( D => n5414, CP => CLK_I, Q => 
                           n_2015, QN => n505);
   KEY_EXPAN0_reg_55_12_inst : FD1 port map( D => n5413, CP => CLK_I, Q => 
                           n_2016, QN => n1583);
   KEY_EXPAN0_reg_54_12_inst : FD1 port map( D => n5412, CP => CLK_I, Q => 
                           n_2017, QN => n512);
   KEY_EXPAN0_reg_53_12_inst : FD1 port map( D => n5411, CP => CLK_I, Q => 
                           n_2018, QN => n1582);
   KEY_EXPAN0_reg_52_12_inst : FD1 port map( D => n5410, CP => CLK_I, Q => 
                           n_2019, QN => n511);
   KEY_EXPAN0_reg_51_12_inst : FD1 port map( D => n5409, CP => CLK_I, Q => 
                           n_2020, QN => n1581);
   KEY_EXPAN0_reg_50_12_inst : FD1 port map( D => n5408, CP => CLK_I, Q => 
                           n_2021, QN => n510);
   KEY_EXPAN0_reg_49_12_inst : FD1 port map( D => n5407, CP => CLK_I, Q => 
                           n_2022, QN => n1580);
   KEY_EXPAN0_reg_48_12_inst : FD1 port map( D => n5406, CP => CLK_I, Q => 
                           n_2023, QN => n509);
   KEY_EXPAN0_reg_47_12_inst : FD1 port map( D => n5405, CP => CLK_I, Q => 
                           n_2024, QN => n1587);
   KEY_EXPAN0_reg_46_12_inst : FD1 port map( D => n5404, CP => CLK_I, Q => 
                           n_2025, QN => n516);
   KEY_EXPAN0_reg_45_12_inst : FD1 port map( D => n5403, CP => CLK_I, Q => 
                           n_2026, QN => n1586);
   KEY_EXPAN0_reg_44_12_inst : FD1 port map( D => n5402, CP => CLK_I, Q => 
                           n_2027, QN => n515);
   KEY_EXPAN0_reg_43_12_inst : FD1 port map( D => n5401, CP => CLK_I, Q => 
                           n_2028, QN => n1585);
   KEY_EXPAN0_reg_42_12_inst : FD1 port map( D => n5400, CP => CLK_I, Q => 
                           n_2029, QN => n514);
   KEY_EXPAN0_reg_41_12_inst : FD1 port map( D => n5399, CP => CLK_I, Q => 
                           n_2030, QN => n1584);
   KEY_EXPAN0_reg_40_12_inst : FD1 port map( D => n5398, CP => CLK_I, Q => 
                           n_2031, QN => n513);
   KEY_EXPAN0_reg_39_12_inst : FD1 port map( D => n5397, CP => CLK_I, Q => 
                           n_2032, QN => n1591);
   KEY_EXPAN0_reg_38_12_inst : FD1 port map( D => n5396, CP => CLK_I, Q => 
                           n_2033, QN => n520);
   KEY_EXPAN0_reg_37_12_inst : FD1 port map( D => n5395, CP => CLK_I, Q => 
                           n_2034, QN => n1590);
   KEY_EXPAN0_reg_36_12_inst : FD1 port map( D => n5394, CP => CLK_I, Q => 
                           n_2035, QN => n519);
   KEY_EXPAN0_reg_35_12_inst : FD1 port map( D => n5393, CP => CLK_I, Q => 
                           n_2036, QN => n1589);
   KEY_EXPAN0_reg_34_12_inst : FD1 port map( D => n5392, CP => CLK_I, Q => 
                           n_2037, QN => n518);
   KEY_EXPAN0_reg_33_12_inst : FD1 port map( D => n5391, CP => CLK_I, Q => 
                           n_2038, QN => n1588);
   KEY_EXPAN0_reg_32_12_inst : FD1 port map( D => n5390, CP => CLK_I, Q => 
                           n_2039, QN => n517);
   KEY_EXPAN0_reg_31_12_inst : FD1 port map( D => n5389, CP => CLK_I, Q => 
                           n_2040, QN => n1563);
   KEY_EXPAN0_reg_30_12_inst : FD1 port map( D => n5388, CP => CLK_I, Q => 
                           n_2041, QN => n492);
   KEY_EXPAN0_reg_29_12_inst : FD1 port map( D => n5387, CP => CLK_I, Q => 
                           n_2042, QN => n1562);
   KEY_EXPAN0_reg_28_12_inst : FD1 port map( D => n5386, CP => CLK_I, Q => 
                           n_2043, QN => n491);
   KEY_EXPAN0_reg_27_12_inst : FD1 port map( D => n5385, CP => CLK_I, Q => 
                           n_2044, QN => n1561);
   KEY_EXPAN0_reg_26_12_inst : FD1 port map( D => n5384, CP => CLK_I, Q => 
                           n_2045, QN => n490);
   KEY_EXPAN0_reg_25_12_inst : FD1 port map( D => n5383, CP => CLK_I, Q => 
                           n_2046, QN => n1560);
   KEY_EXPAN0_reg_24_12_inst : FD1 port map( D => n5382, CP => CLK_I, Q => 
                           n_2047, QN => n489);
   KEY_EXPAN0_reg_23_12_inst : FD1 port map( D => n5381, CP => CLK_I, Q => 
                           n_2048, QN => n1567);
   KEY_EXPAN0_reg_22_12_inst : FD1 port map( D => n5380, CP => CLK_I, Q => 
                           n_2049, QN => n496);
   KEY_EXPAN0_reg_21_12_inst : FD1 port map( D => n5379, CP => CLK_I, Q => 
                           n_2050, QN => n1566);
   KEY_EXPAN0_reg_20_12_inst : FD1 port map( D => n5378, CP => CLK_I, Q => 
                           n_2051, QN => n495);
   KEY_EXPAN0_reg_19_12_inst : FD1 port map( D => n5377, CP => CLK_I, Q => 
                           n_2052, QN => n1565);
   KEY_EXPAN0_reg_18_12_inst : FD1 port map( D => n5376, CP => CLK_I, Q => 
                           n_2053, QN => n494);
   KEY_EXPAN0_reg_17_12_inst : FD1 port map( D => n5375, CP => CLK_I, Q => 
                           n_2054, QN => n1564);
   KEY_EXPAN0_reg_16_12_inst : FD1 port map( D => n5374, CP => CLK_I, Q => 
                           n_2055, QN => n493);
   KEY_EXPAN0_reg_15_12_inst : FD1 port map( D => n5373, CP => CLK_I, Q => 
                           n_2056, QN => n1571);
   KEY_EXPAN0_reg_14_12_inst : FD1 port map( D => n5372, CP => CLK_I, Q => 
                           n_2057, QN => n500);
   KEY_EXPAN0_reg_13_12_inst : FD1 port map( D => n5371, CP => CLK_I, Q => 
                           n_2058, QN => n1570);
   KEY_EXPAN0_reg_12_12_inst : FD1 port map( D => n5370, CP => CLK_I, Q => 
                           n_2059, QN => n499);
   KEY_EXPAN0_reg_11_12_inst : FD1 port map( D => n5369, CP => CLK_I, Q => 
                           n_2060, QN => n1569);
   KEY_EXPAN0_reg_10_12_inst : FD1 port map( D => n5368, CP => CLK_I, Q => 
                           n_2061, QN => n498);
   KEY_EXPAN0_reg_9_12_inst : FD1 port map( D => n5367, CP => CLK_I, Q => 
                           n_2062, QN => n1568);
   KEY_EXPAN0_reg_8_12_inst : FD1 port map( D => n5366, CP => CLK_I, Q => 
                           n_2063, QN => n497);
   KEY_EXPAN0_reg_7_12_inst : FD1 port map( D => n5365, CP => CLK_I, Q => 
                           n_2064, QN => n1575);
   KEY_EXPAN0_reg_6_12_inst : FD1 port map( D => n5364, CP => CLK_I, Q => 
                           n_2065, QN => n504);
   KEY_EXPAN0_reg_5_12_inst : FD1 port map( D => n5363, CP => CLK_I, Q => 
                           n_2066, QN => n1574);
   KEY_EXPAN0_reg_4_12_inst : FD1 port map( D => n5362, CP => CLK_I, Q => 
                           n_2067, QN => n503);
   KEY_EXPAN0_reg_3_12_inst : FD1 port map( D => n5361, CP => CLK_I, Q => 
                           n_2068, QN => n1573);
   KEY_EXPAN0_reg_2_12_inst : FD1 port map( D => n5360, CP => CLK_I, Q => 
                           n_2069, QN => n502);
   KEY_EXPAN0_reg_1_12_inst : FD1 port map( D => n5359, CP => CLK_I, Q => 
                           n_2070, QN => n1572);
   KEY_EXPAN0_reg_0_12_inst : FD1 port map( D => n5358, CP => CLK_I, Q => 
                           n_2071, QN => n501);
   v_KEY_COL_OUT0_reg_12_inst : FD1 port map( D => n4565, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_12_port, QN => n1071);
   v_TEMP_VECTOR_reg_3_inst : FD1 port map( D => n6692, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_3_port, QN => n_2072);
   KEY_EXPAN0_reg_63_3_inst : FD1 port map( D => n4845, CP => CLK_I, Q => 
                           n_2073, QN => n1611);
   KEY_EXPAN0_reg_62_3_inst : FD1 port map( D => n4844, CP => CLK_I, Q => 
                           n_2074, QN => n540);
   KEY_EXPAN0_reg_61_3_inst : FD1 port map( D => n4843, CP => CLK_I, Q => 
                           n_2075, QN => n1610);
   KEY_EXPAN0_reg_60_3_inst : FD1 port map( D => n4842, CP => CLK_I, Q => 
                           n_2076, QN => n539);
   KEY_EXPAN0_reg_59_3_inst : FD1 port map( D => n4841, CP => CLK_I, Q => 
                           n_2077, QN => n1609);
   KEY_EXPAN0_reg_58_3_inst : FD1 port map( D => n4840, CP => CLK_I, Q => 
                           n_2078, QN => n538);
   KEY_EXPAN0_reg_57_3_inst : FD1 port map( D => n4839, CP => CLK_I, Q => 
                           n_2079, QN => n1608);
   KEY_EXPAN0_reg_56_3_inst : FD1 port map( D => n4838, CP => CLK_I, Q => 
                           n_2080, QN => n537);
   KEY_EXPAN0_reg_55_3_inst : FD1 port map( D => n4837, CP => CLK_I, Q => 
                           n_2081, QN => n1615);
   KEY_EXPAN0_reg_54_3_inst : FD1 port map( D => n4836, CP => CLK_I, Q => 
                           n_2082, QN => n544);
   KEY_EXPAN0_reg_53_3_inst : FD1 port map( D => n4835, CP => CLK_I, Q => 
                           n_2083, QN => n1614);
   KEY_EXPAN0_reg_52_3_inst : FD1 port map( D => n4834, CP => CLK_I, Q => 
                           n_2084, QN => n543);
   KEY_EXPAN0_reg_51_3_inst : FD1 port map( D => n4833, CP => CLK_I, Q => 
                           n_2085, QN => n1613);
   KEY_EXPAN0_reg_50_3_inst : FD1 port map( D => n4832, CP => CLK_I, Q => 
                           n_2086, QN => n542);
   KEY_EXPAN0_reg_49_3_inst : FD1 port map( D => n4831, CP => CLK_I, Q => 
                           n_2087, QN => n1612);
   KEY_EXPAN0_reg_48_3_inst : FD1 port map( D => n4830, CP => CLK_I, Q => 
                           n_2088, QN => n541);
   KEY_EXPAN0_reg_47_3_inst : FD1 port map( D => n4829, CP => CLK_I, Q => 
                           n_2089, QN => n1619);
   KEY_EXPAN0_reg_46_3_inst : FD1 port map( D => n4828, CP => CLK_I, Q => 
                           n_2090, QN => n548);
   KEY_EXPAN0_reg_45_3_inst : FD1 port map( D => n4827, CP => CLK_I, Q => 
                           n_2091, QN => n1618);
   KEY_EXPAN0_reg_44_3_inst : FD1 port map( D => n4826, CP => CLK_I, Q => 
                           n_2092, QN => n547);
   KEY_EXPAN0_reg_43_3_inst : FD1 port map( D => n4825, CP => CLK_I, Q => 
                           n_2093, QN => n1617);
   KEY_EXPAN0_reg_42_3_inst : FD1 port map( D => n4824, CP => CLK_I, Q => 
                           n_2094, QN => n546);
   KEY_EXPAN0_reg_41_3_inst : FD1 port map( D => n4823, CP => CLK_I, Q => 
                           n_2095, QN => n1616);
   KEY_EXPAN0_reg_40_3_inst : FD1 port map( D => n4822, CP => CLK_I, Q => 
                           n_2096, QN => n545);
   KEY_EXPAN0_reg_39_3_inst : FD1 port map( D => n4821, CP => CLK_I, Q => 
                           n_2097, QN => n1623);
   KEY_EXPAN0_reg_38_3_inst : FD1 port map( D => n4820, CP => CLK_I, Q => 
                           n_2098, QN => n552);
   KEY_EXPAN0_reg_37_3_inst : FD1 port map( D => n4819, CP => CLK_I, Q => 
                           n_2099, QN => n1622);
   KEY_EXPAN0_reg_36_3_inst : FD1 port map( D => n4818, CP => CLK_I, Q => 
                           n_2100, QN => n551);
   KEY_EXPAN0_reg_35_3_inst : FD1 port map( D => n4817, CP => CLK_I, Q => 
                           n_2101, QN => n1621);
   KEY_EXPAN0_reg_34_3_inst : FD1 port map( D => n4816, CP => CLK_I, Q => 
                           n_2102, QN => n550);
   KEY_EXPAN0_reg_33_3_inst : FD1 port map( D => n4815, CP => CLK_I, Q => 
                           n_2103, QN => n1620);
   KEY_EXPAN0_reg_32_3_inst : FD1 port map( D => n4814, CP => CLK_I, Q => 
                           n_2104, QN => n549);
   KEY_EXPAN0_reg_31_3_inst : FD1 port map( D => n4813, CP => CLK_I, Q => 
                           n_2105, QN => n1595);
   KEY_EXPAN0_reg_30_3_inst : FD1 port map( D => n4812, CP => CLK_I, Q => 
                           n_2106, QN => n524);
   KEY_EXPAN0_reg_29_3_inst : FD1 port map( D => n4811, CP => CLK_I, Q => 
                           n_2107, QN => n1594);
   KEY_EXPAN0_reg_28_3_inst : FD1 port map( D => n4810, CP => CLK_I, Q => 
                           n_2108, QN => n523);
   KEY_EXPAN0_reg_27_3_inst : FD1 port map( D => n4809, CP => CLK_I, Q => 
                           n_2109, QN => n1593);
   KEY_EXPAN0_reg_26_3_inst : FD1 port map( D => n4808, CP => CLK_I, Q => 
                           n_2110, QN => n522);
   KEY_EXPAN0_reg_25_3_inst : FD1 port map( D => n4807, CP => CLK_I, Q => 
                           n_2111, QN => n1592);
   KEY_EXPAN0_reg_24_3_inst : FD1 port map( D => n4806, CP => CLK_I, Q => 
                           n_2112, QN => n521);
   KEY_EXPAN0_reg_23_3_inst : FD1 port map( D => n4805, CP => CLK_I, Q => 
                           n_2113, QN => n1599);
   KEY_EXPAN0_reg_22_3_inst : FD1 port map( D => n4804, CP => CLK_I, Q => 
                           n_2114, QN => n528);
   KEY_EXPAN0_reg_21_3_inst : FD1 port map( D => n4803, CP => CLK_I, Q => 
                           n_2115, QN => n1598);
   KEY_EXPAN0_reg_20_3_inst : FD1 port map( D => n4802, CP => CLK_I, Q => 
                           n_2116, QN => n527);
   KEY_EXPAN0_reg_19_3_inst : FD1 port map( D => n4801, CP => CLK_I, Q => 
                           n_2117, QN => n1597);
   KEY_EXPAN0_reg_18_3_inst : FD1 port map( D => n4800, CP => CLK_I, Q => 
                           n_2118, QN => n526);
   KEY_EXPAN0_reg_17_3_inst : FD1 port map( D => n4799, CP => CLK_I, Q => 
                           n_2119, QN => n1596);
   KEY_EXPAN0_reg_16_3_inst : FD1 port map( D => n4798, CP => CLK_I, Q => 
                           n_2120, QN => n525);
   KEY_EXPAN0_reg_15_3_inst : FD1 port map( D => n4797, CP => CLK_I, Q => 
                           n_2121, QN => n1603);
   KEY_EXPAN0_reg_14_3_inst : FD1 port map( D => n4796, CP => CLK_I, Q => 
                           n_2122, QN => n532);
   KEY_EXPAN0_reg_13_3_inst : FD1 port map( D => n4795, CP => CLK_I, Q => 
                           n_2123, QN => n1602);
   KEY_EXPAN0_reg_12_3_inst : FD1 port map( D => n4794, CP => CLK_I, Q => 
                           n_2124, QN => n531);
   KEY_EXPAN0_reg_11_3_inst : FD1 port map( D => n4793, CP => CLK_I, Q => 
                           n_2125, QN => n1601);
   KEY_EXPAN0_reg_10_3_inst : FD1 port map( D => n4792, CP => CLK_I, Q => 
                           n_2126, QN => n530);
   KEY_EXPAN0_reg_9_3_inst : FD1 port map( D => n4791, CP => CLK_I, Q => n_2127
                           , QN => n1600);
   KEY_EXPAN0_reg_8_3_inst : FD1 port map( D => n4790, CP => CLK_I, Q => n_2128
                           , QN => n529);
   KEY_EXPAN0_reg_7_3_inst : FD1 port map( D => n4789, CP => CLK_I, Q => n_2129
                           , QN => n1607);
   KEY_EXPAN0_reg_6_3_inst : FD1 port map( D => n4788, CP => CLK_I, Q => n_2130
                           , QN => n536);
   KEY_EXPAN0_reg_5_3_inst : FD1 port map( D => n4787, CP => CLK_I, Q => n_2131
                           , QN => n1606);
   KEY_EXPAN0_reg_4_3_inst : FD1 port map( D => n4786, CP => CLK_I, Q => n_2132
                           , QN => n535);
   KEY_EXPAN0_reg_3_3_inst : FD1 port map( D => n4785, CP => CLK_I, Q => n_2133
                           , QN => n1605);
   KEY_EXPAN0_reg_2_3_inst : FD1 port map( D => n4784, CP => CLK_I, Q => n_2134
                           , QN => n534);
   KEY_EXPAN0_reg_1_3_inst : FD1 port map( D => n4783, CP => CLK_I, Q => n_2135
                           , QN => n1604);
   KEY_EXPAN0_reg_0_3_inst : FD1 port map( D => n4782, CP => CLK_I, Q => n_2136
                           , QN => n533);
   v_KEY_COL_OUT0_reg_3_inst : FD1 port map( D => n4564, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_3_port, QN => n1049);
   v_TEMP_VECTOR_reg_27_inst : FD1 port map( D => n6668, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_27_port, QN => n_2137);
   KEY_EXPAN0_reg_63_27_inst : FD1 port map( D => n6381, CP => CLK_I, Q => 
                           n_2138, QN => n1643);
   KEY_EXPAN0_reg_62_27_inst : FD1 port map( D => n6380, CP => CLK_I, Q => 
                           n_2139, QN => n572);
   KEY_EXPAN0_reg_61_27_inst : FD1 port map( D => n6379, CP => CLK_I, Q => 
                           n_2140, QN => n1642);
   KEY_EXPAN0_reg_60_27_inst : FD1 port map( D => n6378, CP => CLK_I, Q => 
                           n_2141, QN => n571);
   KEY_EXPAN0_reg_59_27_inst : FD1 port map( D => n6377, CP => CLK_I, Q => 
                           n_2142, QN => n1641);
   KEY_EXPAN0_reg_58_27_inst : FD1 port map( D => n6376, CP => CLK_I, Q => 
                           n_2143, QN => n570);
   KEY_EXPAN0_reg_57_27_inst : FD1 port map( D => n6375, CP => CLK_I, Q => 
                           n_2144, QN => n1640);
   KEY_EXPAN0_reg_56_27_inst : FD1 port map( D => n6374, CP => CLK_I, Q => 
                           n_2145, QN => n569);
   KEY_EXPAN0_reg_55_27_inst : FD1 port map( D => n6373, CP => CLK_I, Q => 
                           n_2146, QN => n1647);
   KEY_EXPAN0_reg_54_27_inst : FD1 port map( D => n6372, CP => CLK_I, Q => 
                           n_2147, QN => n576);
   KEY_EXPAN0_reg_53_27_inst : FD1 port map( D => n6371, CP => CLK_I, Q => 
                           n_2148, QN => n1646);
   KEY_EXPAN0_reg_52_27_inst : FD1 port map( D => n6370, CP => CLK_I, Q => 
                           n_2149, QN => n575);
   KEY_EXPAN0_reg_51_27_inst : FD1 port map( D => n6369, CP => CLK_I, Q => 
                           n_2150, QN => n1645);
   KEY_EXPAN0_reg_50_27_inst : FD1 port map( D => n6368, CP => CLK_I, Q => 
                           n_2151, QN => n574);
   KEY_EXPAN0_reg_49_27_inst : FD1 port map( D => n6367, CP => CLK_I, Q => 
                           n_2152, QN => n1644);
   KEY_EXPAN0_reg_48_27_inst : FD1 port map( D => n6366, CP => CLK_I, Q => 
                           n_2153, QN => n573);
   KEY_EXPAN0_reg_47_27_inst : FD1 port map( D => n6365, CP => CLK_I, Q => 
                           n_2154, QN => n1651);
   KEY_EXPAN0_reg_46_27_inst : FD1 port map( D => n6364, CP => CLK_I, Q => 
                           n_2155, QN => n580);
   KEY_EXPAN0_reg_45_27_inst : FD1 port map( D => n6363, CP => CLK_I, Q => 
                           n_2156, QN => n1650);
   KEY_EXPAN0_reg_44_27_inst : FD1 port map( D => n6362, CP => CLK_I, Q => 
                           n_2157, QN => n579);
   KEY_EXPAN0_reg_43_27_inst : FD1 port map( D => n6361, CP => CLK_I, Q => 
                           n_2158, QN => n1649);
   KEY_EXPAN0_reg_42_27_inst : FD1 port map( D => n6360, CP => CLK_I, Q => 
                           n_2159, QN => n578);
   KEY_EXPAN0_reg_41_27_inst : FD1 port map( D => n6359, CP => CLK_I, Q => 
                           n_2160, QN => n1648);
   KEY_EXPAN0_reg_40_27_inst : FD1 port map( D => n6358, CP => CLK_I, Q => 
                           n_2161, QN => n577);
   KEY_EXPAN0_reg_39_27_inst : FD1 port map( D => n6357, CP => CLK_I, Q => 
                           n_2162, QN => n1655);
   KEY_EXPAN0_reg_38_27_inst : FD1 port map( D => n6356, CP => CLK_I, Q => 
                           n_2163, QN => n584);
   KEY_EXPAN0_reg_37_27_inst : FD1 port map( D => n6355, CP => CLK_I, Q => 
                           n_2164, QN => n1654);
   KEY_EXPAN0_reg_36_27_inst : FD1 port map( D => n6354, CP => CLK_I, Q => 
                           n_2165, QN => n583);
   KEY_EXPAN0_reg_35_27_inst : FD1 port map( D => n6353, CP => CLK_I, Q => 
                           n_2166, QN => n1653);
   KEY_EXPAN0_reg_34_27_inst : FD1 port map( D => n6352, CP => CLK_I, Q => 
                           n_2167, QN => n582);
   KEY_EXPAN0_reg_33_27_inst : FD1 port map( D => n6351, CP => CLK_I, Q => 
                           n_2168, QN => n1652);
   KEY_EXPAN0_reg_32_27_inst : FD1 port map( D => n6350, CP => CLK_I, Q => 
                           n_2169, QN => n581);
   KEY_EXPAN0_reg_31_27_inst : FD1 port map( D => n6349, CP => CLK_I, Q => 
                           n_2170, QN => n1627);
   KEY_EXPAN0_reg_30_27_inst : FD1 port map( D => n6348, CP => CLK_I, Q => 
                           n_2171, QN => n556);
   KEY_EXPAN0_reg_29_27_inst : FD1 port map( D => n6347, CP => CLK_I, Q => 
                           n_2172, QN => n1626);
   KEY_EXPAN0_reg_28_27_inst : FD1 port map( D => n6346, CP => CLK_I, Q => 
                           n_2173, QN => n555);
   KEY_EXPAN0_reg_27_27_inst : FD1 port map( D => n6345, CP => CLK_I, Q => 
                           n_2174, QN => n1625);
   KEY_EXPAN0_reg_26_27_inst : FD1 port map( D => n6344, CP => CLK_I, Q => 
                           n_2175, QN => n554);
   KEY_EXPAN0_reg_25_27_inst : FD1 port map( D => n6343, CP => CLK_I, Q => 
                           n_2176, QN => n1624);
   KEY_EXPAN0_reg_24_27_inst : FD1 port map( D => n6342, CP => CLK_I, Q => 
                           n_2177, QN => n553);
   KEY_EXPAN0_reg_23_27_inst : FD1 port map( D => n6341, CP => CLK_I, Q => 
                           n_2178, QN => n1631);
   KEY_EXPAN0_reg_22_27_inst : FD1 port map( D => n6340, CP => CLK_I, Q => 
                           n_2179, QN => n560);
   KEY_EXPAN0_reg_21_27_inst : FD1 port map( D => n6339, CP => CLK_I, Q => 
                           n_2180, QN => n1630);
   KEY_EXPAN0_reg_20_27_inst : FD1 port map( D => n6338, CP => CLK_I, Q => 
                           n_2181, QN => n559);
   KEY_EXPAN0_reg_19_27_inst : FD1 port map( D => n6337, CP => CLK_I, Q => 
                           n_2182, QN => n1629);
   KEY_EXPAN0_reg_18_27_inst : FD1 port map( D => n6336, CP => CLK_I, Q => 
                           n_2183, QN => n558);
   KEY_EXPAN0_reg_17_27_inst : FD1 port map( D => n6335, CP => CLK_I, Q => 
                           n_2184, QN => n1628);
   KEY_EXPAN0_reg_16_27_inst : FD1 port map( D => n6334, CP => CLK_I, Q => 
                           n_2185, QN => n557);
   KEY_EXPAN0_reg_15_27_inst : FD1 port map( D => n6333, CP => CLK_I, Q => 
                           n_2186, QN => n1635);
   KEY_EXPAN0_reg_14_27_inst : FD1 port map( D => n6332, CP => CLK_I, Q => 
                           n_2187, QN => n564);
   KEY_EXPAN0_reg_13_27_inst : FD1 port map( D => n6331, CP => CLK_I, Q => 
                           n_2188, QN => n1634);
   KEY_EXPAN0_reg_12_27_inst : FD1 port map( D => n6330, CP => CLK_I, Q => 
                           n_2189, QN => n563);
   KEY_EXPAN0_reg_11_27_inst : FD1 port map( D => n6329, CP => CLK_I, Q => 
                           n_2190, QN => n1633);
   KEY_EXPAN0_reg_10_27_inst : FD1 port map( D => n6328, CP => CLK_I, Q => 
                           n_2191, QN => n562);
   KEY_EXPAN0_reg_9_27_inst : FD1 port map( D => n6327, CP => CLK_I, Q => 
                           n_2192, QN => n1632);
   KEY_EXPAN0_reg_8_27_inst : FD1 port map( D => n6326, CP => CLK_I, Q => 
                           n_2193, QN => n561);
   KEY_EXPAN0_reg_7_27_inst : FD1 port map( D => n6325, CP => CLK_I, Q => 
                           n_2194, QN => n1639);
   KEY_EXPAN0_reg_6_27_inst : FD1 port map( D => n6324, CP => CLK_I, Q => 
                           n_2195, QN => n568);
   KEY_EXPAN0_reg_5_27_inst : FD1 port map( D => n6323, CP => CLK_I, Q => 
                           n_2196, QN => n1638);
   KEY_EXPAN0_reg_4_27_inst : FD1 port map( D => n6322, CP => CLK_I, Q => 
                           n_2197, QN => n567);
   KEY_EXPAN0_reg_3_27_inst : FD1 port map( D => n6321, CP => CLK_I, Q => 
                           n_2198, QN => n1637);
   KEY_EXPAN0_reg_2_27_inst : FD1 port map( D => n6320, CP => CLK_I, Q => 
                           n_2199, QN => n566);
   KEY_EXPAN0_reg_1_27_inst : FD1 port map( D => n6319, CP => CLK_I, Q => 
                           n_2200, QN => n1636);
   KEY_EXPAN0_reg_0_27_inst : FD1 port map( D => n6318, CP => CLK_I, Q => 
                           n_2201, QN => n565);
   v_KEY_COL_OUT0_reg_27_inst : FD1 port map( D => n4563, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_27_port, QN => n1055);
   v_TEMP_VECTOR_reg_19_inst : FD1 port map( D => n6676, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_19_port, QN => n_2202);
   KEY_EXPAN0_reg_63_19_inst : FD1 port map( D => n5869, CP => CLK_I, Q => 
                           n_2203, QN => n1675);
   KEY_EXPAN0_reg_62_19_inst : FD1 port map( D => n5868, CP => CLK_I, Q => 
                           n_2204, QN => n604);
   KEY_EXPAN0_reg_61_19_inst : FD1 port map( D => n5867, CP => CLK_I, Q => 
                           n_2205, QN => n1674);
   KEY_EXPAN0_reg_60_19_inst : FD1 port map( D => n5866, CP => CLK_I, Q => 
                           n_2206, QN => n603);
   KEY_EXPAN0_reg_59_19_inst : FD1 port map( D => n5865, CP => CLK_I, Q => 
                           n_2207, QN => n1673);
   KEY_EXPAN0_reg_58_19_inst : FD1 port map( D => n5864, CP => CLK_I, Q => 
                           n_2208, QN => n602);
   KEY_EXPAN0_reg_57_19_inst : FD1 port map( D => n5863, CP => CLK_I, Q => 
                           n_2209, QN => n1672);
   KEY_EXPAN0_reg_56_19_inst : FD1 port map( D => n5862, CP => CLK_I, Q => 
                           n_2210, QN => n601);
   KEY_EXPAN0_reg_55_19_inst : FD1 port map( D => n5861, CP => CLK_I, Q => 
                           n_2211, QN => n1679);
   KEY_EXPAN0_reg_54_19_inst : FD1 port map( D => n5860, CP => CLK_I, Q => 
                           n_2212, QN => n608);
   KEY_EXPAN0_reg_53_19_inst : FD1 port map( D => n5859, CP => CLK_I, Q => 
                           n_2213, QN => n1678);
   KEY_EXPAN0_reg_52_19_inst : FD1 port map( D => n5858, CP => CLK_I, Q => 
                           n_2214, QN => n607);
   KEY_EXPAN0_reg_51_19_inst : FD1 port map( D => n5857, CP => CLK_I, Q => 
                           n_2215, QN => n1677);
   KEY_EXPAN0_reg_50_19_inst : FD1 port map( D => n5856, CP => CLK_I, Q => 
                           n_2216, QN => n606);
   KEY_EXPAN0_reg_49_19_inst : FD1 port map( D => n5855, CP => CLK_I, Q => 
                           n_2217, QN => n1676);
   KEY_EXPAN0_reg_48_19_inst : FD1 port map( D => n5854, CP => CLK_I, Q => 
                           n_2218, QN => n605);
   KEY_EXPAN0_reg_47_19_inst : FD1 port map( D => n5853, CP => CLK_I, Q => 
                           n_2219, QN => n1683);
   KEY_EXPAN0_reg_46_19_inst : FD1 port map( D => n5852, CP => CLK_I, Q => 
                           n_2220, QN => n612);
   KEY_EXPAN0_reg_45_19_inst : FD1 port map( D => n5851, CP => CLK_I, Q => 
                           n_2221, QN => n1682);
   KEY_EXPAN0_reg_44_19_inst : FD1 port map( D => n5850, CP => CLK_I, Q => 
                           n_2222, QN => n611);
   KEY_EXPAN0_reg_43_19_inst : FD1 port map( D => n5849, CP => CLK_I, Q => 
                           n_2223, QN => n1681);
   KEY_EXPAN0_reg_42_19_inst : FD1 port map( D => n5848, CP => CLK_I, Q => 
                           n_2224, QN => n610);
   KEY_EXPAN0_reg_41_19_inst : FD1 port map( D => n5847, CP => CLK_I, Q => 
                           n_2225, QN => n1680);
   KEY_EXPAN0_reg_40_19_inst : FD1 port map( D => n5846, CP => CLK_I, Q => 
                           n_2226, QN => n609);
   KEY_EXPAN0_reg_39_19_inst : FD1 port map( D => n5845, CP => CLK_I, Q => 
                           n_2227, QN => n1687);
   KEY_EXPAN0_reg_38_19_inst : FD1 port map( D => n5844, CP => CLK_I, Q => 
                           n_2228, QN => n616);
   KEY_EXPAN0_reg_37_19_inst : FD1 port map( D => n5843, CP => CLK_I, Q => 
                           n_2229, QN => n1686);
   KEY_EXPAN0_reg_36_19_inst : FD1 port map( D => n5842, CP => CLK_I, Q => 
                           n_2230, QN => n615);
   KEY_EXPAN0_reg_35_19_inst : FD1 port map( D => n5841, CP => CLK_I, Q => 
                           n_2231, QN => n1685);
   KEY_EXPAN0_reg_34_19_inst : FD1 port map( D => n5840, CP => CLK_I, Q => 
                           n_2232, QN => n614);
   KEY_EXPAN0_reg_33_19_inst : FD1 port map( D => n5839, CP => CLK_I, Q => 
                           n_2233, QN => n1684);
   KEY_EXPAN0_reg_32_19_inst : FD1 port map( D => n5838, CP => CLK_I, Q => 
                           n_2234, QN => n613);
   KEY_EXPAN0_reg_31_19_inst : FD1 port map( D => n5837, CP => CLK_I, Q => 
                           n_2235, QN => n1659);
   KEY_EXPAN0_reg_30_19_inst : FD1 port map( D => n5836, CP => CLK_I, Q => 
                           n_2236, QN => n588);
   KEY_EXPAN0_reg_29_19_inst : FD1 port map( D => n5835, CP => CLK_I, Q => 
                           n_2237, QN => n1658);
   KEY_EXPAN0_reg_28_19_inst : FD1 port map( D => n5834, CP => CLK_I, Q => 
                           n_2238, QN => n587);
   KEY_EXPAN0_reg_27_19_inst : FD1 port map( D => n5833, CP => CLK_I, Q => 
                           n_2239, QN => n1657);
   KEY_EXPAN0_reg_26_19_inst : FD1 port map( D => n5832, CP => CLK_I, Q => 
                           n_2240, QN => n586);
   KEY_EXPAN0_reg_25_19_inst : FD1 port map( D => n5831, CP => CLK_I, Q => 
                           n_2241, QN => n1656);
   KEY_EXPAN0_reg_24_19_inst : FD1 port map( D => n5830, CP => CLK_I, Q => 
                           n_2242, QN => n585);
   KEY_EXPAN0_reg_23_19_inst : FD1 port map( D => n5829, CP => CLK_I, Q => 
                           n_2243, QN => n1663);
   KEY_EXPAN0_reg_22_19_inst : FD1 port map( D => n5828, CP => CLK_I, Q => 
                           n_2244, QN => n592);
   KEY_EXPAN0_reg_21_19_inst : FD1 port map( D => n5827, CP => CLK_I, Q => 
                           n_2245, QN => n1662);
   KEY_EXPAN0_reg_20_19_inst : FD1 port map( D => n5826, CP => CLK_I, Q => 
                           n_2246, QN => n591);
   KEY_EXPAN0_reg_19_19_inst : FD1 port map( D => n5825, CP => CLK_I, Q => 
                           n_2247, QN => n1661);
   KEY_EXPAN0_reg_18_19_inst : FD1 port map( D => n5824, CP => CLK_I, Q => 
                           n_2248, QN => n590);
   KEY_EXPAN0_reg_17_19_inst : FD1 port map( D => n5823, CP => CLK_I, Q => 
                           n_2249, QN => n1660);
   KEY_EXPAN0_reg_16_19_inst : FD1 port map( D => n5822, CP => CLK_I, Q => 
                           n_2250, QN => n589);
   KEY_EXPAN0_reg_15_19_inst : FD1 port map( D => n5821, CP => CLK_I, Q => 
                           n_2251, QN => n1667);
   KEY_EXPAN0_reg_14_19_inst : FD1 port map( D => n5820, CP => CLK_I, Q => 
                           n_2252, QN => n596);
   KEY_EXPAN0_reg_13_19_inst : FD1 port map( D => n5819, CP => CLK_I, Q => 
                           n_2253, QN => n1666);
   KEY_EXPAN0_reg_12_19_inst : FD1 port map( D => n5818, CP => CLK_I, Q => 
                           n_2254, QN => n595);
   KEY_EXPAN0_reg_11_19_inst : FD1 port map( D => n5817, CP => CLK_I, Q => 
                           n_2255, QN => n1665);
   KEY_EXPAN0_reg_10_19_inst : FD1 port map( D => n5816, CP => CLK_I, Q => 
                           n_2256, QN => n594);
   KEY_EXPAN0_reg_9_19_inst : FD1 port map( D => n5815, CP => CLK_I, Q => 
                           n_2257, QN => n1664);
   KEY_EXPAN0_reg_8_19_inst : FD1 port map( D => n5814, CP => CLK_I, Q => 
                           n_2258, QN => n593);
   KEY_EXPAN0_reg_7_19_inst : FD1 port map( D => n5813, CP => CLK_I, Q => 
                           n_2259, QN => n1671);
   KEY_EXPAN0_reg_6_19_inst : FD1 port map( D => n5812, CP => CLK_I, Q => 
                           n_2260, QN => n600);
   KEY_EXPAN0_reg_5_19_inst : FD1 port map( D => n5811, CP => CLK_I, Q => 
                           n_2261, QN => n1670);
   KEY_EXPAN0_reg_4_19_inst : FD1 port map( D => n5810, CP => CLK_I, Q => 
                           n_2262, QN => n599);
   KEY_EXPAN0_reg_3_19_inst : FD1 port map( D => n5809, CP => CLK_I, Q => 
                           n_2263, QN => n1669);
   KEY_EXPAN0_reg_2_19_inst : FD1 port map( D => n5808, CP => CLK_I, Q => 
                           n_2264, QN => n598);
   KEY_EXPAN0_reg_1_19_inst : FD1 port map( D => n5807, CP => CLK_I, Q => 
                           n_2265, QN => n1668);
   KEY_EXPAN0_reg_0_19_inst : FD1 port map( D => n5806, CP => CLK_I, Q => 
                           n_2266, QN => n597);
   v_KEY_COL_OUT0_reg_19_inst : FD1 port map( D => n4562, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_19_port, QN => n1064);
   v_TEMP_VECTOR_reg_11_inst : FD1 port map( D => n6684, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_11_port, QN => n_2267);
   KEY_EXPAN0_reg_63_11_inst : FD1 port map( D => n5357, CP => CLK_I, Q => 
                           n_2268, QN => n1707);
   KEY_EXPAN0_reg_62_11_inst : FD1 port map( D => n5356, CP => CLK_I, Q => 
                           n_2269, QN => n636);
   KEY_EXPAN0_reg_61_11_inst : FD1 port map( D => n5355, CP => CLK_I, Q => 
                           n_2270, QN => n1706);
   KEY_EXPAN0_reg_60_11_inst : FD1 port map( D => n5354, CP => CLK_I, Q => 
                           n_2271, QN => n635);
   KEY_EXPAN0_reg_59_11_inst : FD1 port map( D => n5353, CP => CLK_I, Q => 
                           n_2272, QN => n1705);
   KEY_EXPAN0_reg_58_11_inst : FD1 port map( D => n5352, CP => CLK_I, Q => 
                           n_2273, QN => n634);
   KEY_EXPAN0_reg_57_11_inst : FD1 port map( D => n5351, CP => CLK_I, Q => 
                           n_2274, QN => n1704);
   KEY_EXPAN0_reg_56_11_inst : FD1 port map( D => n5350, CP => CLK_I, Q => 
                           n_2275, QN => n633);
   KEY_EXPAN0_reg_55_11_inst : FD1 port map( D => n5349, CP => CLK_I, Q => 
                           n_2276, QN => n1711);
   KEY_EXPAN0_reg_54_11_inst : FD1 port map( D => n5348, CP => CLK_I, Q => 
                           n_2277, QN => n640);
   KEY_EXPAN0_reg_53_11_inst : FD1 port map( D => n5347, CP => CLK_I, Q => 
                           n_2278, QN => n1710);
   KEY_EXPAN0_reg_52_11_inst : FD1 port map( D => n5346, CP => CLK_I, Q => 
                           n_2279, QN => n639);
   KEY_EXPAN0_reg_51_11_inst : FD1 port map( D => n5345, CP => CLK_I, Q => 
                           n_2280, QN => n1709);
   KEY_EXPAN0_reg_50_11_inst : FD1 port map( D => n5344, CP => CLK_I, Q => 
                           n_2281, QN => n638);
   KEY_EXPAN0_reg_49_11_inst : FD1 port map( D => n5343, CP => CLK_I, Q => 
                           n_2282, QN => n1708);
   KEY_EXPAN0_reg_48_11_inst : FD1 port map( D => n5342, CP => CLK_I, Q => 
                           n_2283, QN => n637);
   KEY_EXPAN0_reg_47_11_inst : FD1 port map( D => n5341, CP => CLK_I, Q => 
                           n_2284, QN => n1715);
   KEY_EXPAN0_reg_46_11_inst : FD1 port map( D => n5340, CP => CLK_I, Q => 
                           n_2285, QN => n644);
   KEY_EXPAN0_reg_45_11_inst : FD1 port map( D => n5339, CP => CLK_I, Q => 
                           n_2286, QN => n1714);
   KEY_EXPAN0_reg_44_11_inst : FD1 port map( D => n5338, CP => CLK_I, Q => 
                           n_2287, QN => n643);
   KEY_EXPAN0_reg_43_11_inst : FD1 port map( D => n5337, CP => CLK_I, Q => 
                           n_2288, QN => n1713);
   KEY_EXPAN0_reg_42_11_inst : FD1 port map( D => n5336, CP => CLK_I, Q => 
                           n_2289, QN => n642);
   KEY_EXPAN0_reg_41_11_inst : FD1 port map( D => n5335, CP => CLK_I, Q => 
                           n_2290, QN => n1712);
   KEY_EXPAN0_reg_40_11_inst : FD1 port map( D => n5334, CP => CLK_I, Q => 
                           n_2291, QN => n641);
   KEY_EXPAN0_reg_39_11_inst : FD1 port map( D => n5333, CP => CLK_I, Q => 
                           n_2292, QN => n1719);
   KEY_EXPAN0_reg_38_11_inst : FD1 port map( D => n5332, CP => CLK_I, Q => 
                           n_2293, QN => n648);
   KEY_EXPAN0_reg_37_11_inst : FD1 port map( D => n5331, CP => CLK_I, Q => 
                           n_2294, QN => n1718);
   KEY_EXPAN0_reg_36_11_inst : FD1 port map( D => n5330, CP => CLK_I, Q => 
                           n_2295, QN => n647);
   KEY_EXPAN0_reg_35_11_inst : FD1 port map( D => n5329, CP => CLK_I, Q => 
                           n_2296, QN => n1717);
   KEY_EXPAN0_reg_34_11_inst : FD1 port map( D => n5328, CP => CLK_I, Q => 
                           n_2297, QN => n646);
   KEY_EXPAN0_reg_33_11_inst : FD1 port map( D => n5327, CP => CLK_I, Q => 
                           n_2298, QN => n1716);
   KEY_EXPAN0_reg_32_11_inst : FD1 port map( D => n5326, CP => CLK_I, Q => 
                           n_2299, QN => n645);
   KEY_EXPAN0_reg_31_11_inst : FD1 port map( D => n5325, CP => CLK_I, Q => 
                           n_2300, QN => n1691);
   KEY_EXPAN0_reg_30_11_inst : FD1 port map( D => n5324, CP => CLK_I, Q => 
                           n_2301, QN => n620);
   KEY_EXPAN0_reg_29_11_inst : FD1 port map( D => n5323, CP => CLK_I, Q => 
                           n_2302, QN => n1690);
   KEY_EXPAN0_reg_28_11_inst : FD1 port map( D => n5322, CP => CLK_I, Q => 
                           n_2303, QN => n619);
   KEY_EXPAN0_reg_27_11_inst : FD1 port map( D => n5321, CP => CLK_I, Q => 
                           n_2304, QN => n1689);
   KEY_EXPAN0_reg_26_11_inst : FD1 port map( D => n5320, CP => CLK_I, Q => 
                           n_2305, QN => n618);
   KEY_EXPAN0_reg_25_11_inst : FD1 port map( D => n5319, CP => CLK_I, Q => 
                           n_2306, QN => n1688);
   KEY_EXPAN0_reg_24_11_inst : FD1 port map( D => n5318, CP => CLK_I, Q => 
                           n_2307, QN => n617);
   KEY_EXPAN0_reg_23_11_inst : FD1 port map( D => n5317, CP => CLK_I, Q => 
                           n_2308, QN => n1695);
   KEY_EXPAN0_reg_22_11_inst : FD1 port map( D => n5316, CP => CLK_I, Q => 
                           n_2309, QN => n624);
   KEY_EXPAN0_reg_21_11_inst : FD1 port map( D => n5315, CP => CLK_I, Q => 
                           n_2310, QN => n1694);
   KEY_EXPAN0_reg_20_11_inst : FD1 port map( D => n5314, CP => CLK_I, Q => 
                           n_2311, QN => n623);
   KEY_EXPAN0_reg_19_11_inst : FD1 port map( D => n5313, CP => CLK_I, Q => 
                           n_2312, QN => n1693);
   KEY_EXPAN0_reg_18_11_inst : FD1 port map( D => n5312, CP => CLK_I, Q => 
                           n_2313, QN => n622);
   KEY_EXPAN0_reg_17_11_inst : FD1 port map( D => n5311, CP => CLK_I, Q => 
                           n_2314, QN => n1692);
   KEY_EXPAN0_reg_16_11_inst : FD1 port map( D => n5310, CP => CLK_I, Q => 
                           n_2315, QN => n621);
   KEY_EXPAN0_reg_15_11_inst : FD1 port map( D => n5309, CP => CLK_I, Q => 
                           n_2316, QN => n1699);
   KEY_EXPAN0_reg_14_11_inst : FD1 port map( D => n5308, CP => CLK_I, Q => 
                           n_2317, QN => n628);
   KEY_EXPAN0_reg_13_11_inst : FD1 port map( D => n5307, CP => CLK_I, Q => 
                           n_2318, QN => n1698);
   KEY_EXPAN0_reg_12_11_inst : FD1 port map( D => n5306, CP => CLK_I, Q => 
                           n_2319, QN => n627);
   KEY_EXPAN0_reg_11_11_inst : FD1 port map( D => n5305, CP => CLK_I, Q => 
                           n_2320, QN => n1697);
   KEY_EXPAN0_reg_10_11_inst : FD1 port map( D => n5304, CP => CLK_I, Q => 
                           n_2321, QN => n626);
   KEY_EXPAN0_reg_9_11_inst : FD1 port map( D => n5303, CP => CLK_I, Q => 
                           n_2322, QN => n1696);
   KEY_EXPAN0_reg_8_11_inst : FD1 port map( D => n5302, CP => CLK_I, Q => 
                           n_2323, QN => n625);
   KEY_EXPAN0_reg_7_11_inst : FD1 port map( D => n5301, CP => CLK_I, Q => 
                           n_2324, QN => n1703);
   KEY_EXPAN0_reg_6_11_inst : FD1 port map( D => n5300, CP => CLK_I, Q => 
                           n_2325, QN => n632);
   KEY_EXPAN0_reg_5_11_inst : FD1 port map( D => n5299, CP => CLK_I, Q => 
                           n_2326, QN => n1702);
   KEY_EXPAN0_reg_4_11_inst : FD1 port map( D => n5298, CP => CLK_I, Q => 
                           n_2327, QN => n631);
   KEY_EXPAN0_reg_3_11_inst : FD1 port map( D => n5297, CP => CLK_I, Q => 
                           n_2328, QN => n1701);
   KEY_EXPAN0_reg_2_11_inst : FD1 port map( D => n5296, CP => CLK_I, Q => 
                           n_2329, QN => n630);
   KEY_EXPAN0_reg_1_11_inst : FD1 port map( D => n5295, CP => CLK_I, Q => 
                           n_2330, QN => n1700);
   KEY_EXPAN0_reg_0_11_inst : FD1 port map( D => n5294, CP => CLK_I, Q => 
                           n_2331, QN => n629);
   v_KEY_COL_OUT0_reg_11_inst : FD1 port map( D => n4561, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_11_port, QN => n1072);
   v_TEMP_VECTOR_reg_2_inst : FD1 port map( D => n6693, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_2_port, QN => n_2332);
   KEY_EXPAN0_reg_63_2_inst : FD1 port map( D => n4781, CP => CLK_I, Q => 
                           n_2333, QN => n1739);
   KEY_EXPAN0_reg_62_2_inst : FD1 port map( D => n4780, CP => CLK_I, Q => 
                           n_2334, QN => n668);
   KEY_EXPAN0_reg_61_2_inst : FD1 port map( D => n4779, CP => CLK_I, Q => 
                           n_2335, QN => n1738);
   KEY_EXPAN0_reg_60_2_inst : FD1 port map( D => n4778, CP => CLK_I, Q => 
                           n_2336, QN => n667);
   KEY_EXPAN0_reg_59_2_inst : FD1 port map( D => n4777, CP => CLK_I, Q => 
                           n_2337, QN => n1737);
   KEY_EXPAN0_reg_58_2_inst : FD1 port map( D => n4776, CP => CLK_I, Q => 
                           n_2338, QN => n666);
   KEY_EXPAN0_reg_57_2_inst : FD1 port map( D => n4775, CP => CLK_I, Q => 
                           n_2339, QN => n1736);
   KEY_EXPAN0_reg_56_2_inst : FD1 port map( D => n4774, CP => CLK_I, Q => 
                           n_2340, QN => n665);
   KEY_EXPAN0_reg_55_2_inst : FD1 port map( D => n4773, CP => CLK_I, Q => 
                           n_2341, QN => n1743);
   KEY_EXPAN0_reg_54_2_inst : FD1 port map( D => n4772, CP => CLK_I, Q => 
                           n_2342, QN => n672);
   KEY_EXPAN0_reg_53_2_inst : FD1 port map( D => n4771, CP => CLK_I, Q => 
                           n_2343, QN => n1742);
   KEY_EXPAN0_reg_52_2_inst : FD1 port map( D => n4770, CP => CLK_I, Q => 
                           n_2344, QN => n671);
   KEY_EXPAN0_reg_51_2_inst : FD1 port map( D => n4769, CP => CLK_I, Q => 
                           n_2345, QN => n1741);
   KEY_EXPAN0_reg_50_2_inst : FD1 port map( D => n4768, CP => CLK_I, Q => 
                           n_2346, QN => n670);
   KEY_EXPAN0_reg_49_2_inst : FD1 port map( D => n4767, CP => CLK_I, Q => 
                           n_2347, QN => n1740);
   KEY_EXPAN0_reg_48_2_inst : FD1 port map( D => n4766, CP => CLK_I, Q => 
                           n_2348, QN => n669);
   KEY_EXPAN0_reg_47_2_inst : FD1 port map( D => n4765, CP => CLK_I, Q => 
                           n_2349, QN => n1747);
   KEY_EXPAN0_reg_46_2_inst : FD1 port map( D => n4764, CP => CLK_I, Q => 
                           n_2350, QN => n676);
   KEY_EXPAN0_reg_45_2_inst : FD1 port map( D => n4763, CP => CLK_I, Q => 
                           n_2351, QN => n1746);
   KEY_EXPAN0_reg_44_2_inst : FD1 port map( D => n4762, CP => CLK_I, Q => 
                           n_2352, QN => n675);
   KEY_EXPAN0_reg_43_2_inst : FD1 port map( D => n4761, CP => CLK_I, Q => 
                           n_2353, QN => n1745);
   KEY_EXPAN0_reg_42_2_inst : FD1 port map( D => n4760, CP => CLK_I, Q => 
                           n_2354, QN => n674);
   KEY_EXPAN0_reg_41_2_inst : FD1 port map( D => n4759, CP => CLK_I, Q => 
                           n_2355, QN => n1744);
   KEY_EXPAN0_reg_40_2_inst : FD1 port map( D => n4758, CP => CLK_I, Q => 
                           n_2356, QN => n673);
   KEY_EXPAN0_reg_39_2_inst : FD1 port map( D => n4757, CP => CLK_I, Q => 
                           n_2357, QN => n1751);
   KEY_EXPAN0_reg_38_2_inst : FD1 port map( D => n4756, CP => CLK_I, Q => 
                           n_2358, QN => n680);
   KEY_EXPAN0_reg_37_2_inst : FD1 port map( D => n4755, CP => CLK_I, Q => 
                           n_2359, QN => n1750);
   KEY_EXPAN0_reg_36_2_inst : FD1 port map( D => n4754, CP => CLK_I, Q => 
                           n_2360, QN => n679);
   KEY_EXPAN0_reg_35_2_inst : FD1 port map( D => n4753, CP => CLK_I, Q => 
                           n_2361, QN => n1749);
   KEY_EXPAN0_reg_34_2_inst : FD1 port map( D => n4752, CP => CLK_I, Q => 
                           n_2362, QN => n678);
   KEY_EXPAN0_reg_33_2_inst : FD1 port map( D => n4751, CP => CLK_I, Q => 
                           n_2363, QN => n1748);
   KEY_EXPAN0_reg_32_2_inst : FD1 port map( D => n4750, CP => CLK_I, Q => 
                           n_2364, QN => n677);
   KEY_EXPAN0_reg_31_2_inst : FD1 port map( D => n4749, CP => CLK_I, Q => 
                           n_2365, QN => n1723);
   KEY_EXPAN0_reg_30_2_inst : FD1 port map( D => n4748, CP => CLK_I, Q => 
                           n_2366, QN => n652);
   KEY_EXPAN0_reg_29_2_inst : FD1 port map( D => n4747, CP => CLK_I, Q => 
                           n_2367, QN => n1722);
   KEY_EXPAN0_reg_28_2_inst : FD1 port map( D => n4746, CP => CLK_I, Q => 
                           n_2368, QN => n651);
   KEY_EXPAN0_reg_27_2_inst : FD1 port map( D => n4745, CP => CLK_I, Q => 
                           n_2369, QN => n1721);
   KEY_EXPAN0_reg_26_2_inst : FD1 port map( D => n4744, CP => CLK_I, Q => 
                           n_2370, QN => n650);
   KEY_EXPAN0_reg_25_2_inst : FD1 port map( D => n4743, CP => CLK_I, Q => 
                           n_2371, QN => n1720);
   KEY_EXPAN0_reg_24_2_inst : FD1 port map( D => n4742, CP => CLK_I, Q => 
                           n_2372, QN => n649);
   KEY_EXPAN0_reg_23_2_inst : FD1 port map( D => n4741, CP => CLK_I, Q => 
                           n_2373, QN => n1727);
   KEY_EXPAN0_reg_22_2_inst : FD1 port map( D => n4740, CP => CLK_I, Q => 
                           n_2374, QN => n656);
   KEY_EXPAN0_reg_21_2_inst : FD1 port map( D => n4739, CP => CLK_I, Q => 
                           n_2375, QN => n1726);
   KEY_EXPAN0_reg_20_2_inst : FD1 port map( D => n4738, CP => CLK_I, Q => 
                           n_2376, QN => n655);
   KEY_EXPAN0_reg_19_2_inst : FD1 port map( D => n4737, CP => CLK_I, Q => 
                           n_2377, QN => n1725);
   KEY_EXPAN0_reg_18_2_inst : FD1 port map( D => n4736, CP => CLK_I, Q => 
                           n_2378, QN => n654);
   KEY_EXPAN0_reg_17_2_inst : FD1 port map( D => n4735, CP => CLK_I, Q => 
                           n_2379, QN => n1724);
   KEY_EXPAN0_reg_16_2_inst : FD1 port map( D => n4734, CP => CLK_I, Q => 
                           n_2380, QN => n653);
   KEY_EXPAN0_reg_15_2_inst : FD1 port map( D => n4733, CP => CLK_I, Q => 
                           n_2381, QN => n1731);
   KEY_EXPAN0_reg_14_2_inst : FD1 port map( D => n4732, CP => CLK_I, Q => 
                           n_2382, QN => n660);
   KEY_EXPAN0_reg_13_2_inst : FD1 port map( D => n4731, CP => CLK_I, Q => 
                           n_2383, QN => n1730);
   KEY_EXPAN0_reg_12_2_inst : FD1 port map( D => n4730, CP => CLK_I, Q => 
                           n_2384, QN => n659);
   KEY_EXPAN0_reg_11_2_inst : FD1 port map( D => n4729, CP => CLK_I, Q => 
                           n_2385, QN => n1729);
   KEY_EXPAN0_reg_10_2_inst : FD1 port map( D => n4728, CP => CLK_I, Q => 
                           n_2386, QN => n658);
   KEY_EXPAN0_reg_9_2_inst : FD1 port map( D => n4727, CP => CLK_I, Q => n_2387
                           , QN => n1728);
   KEY_EXPAN0_reg_8_2_inst : FD1 port map( D => n4726, CP => CLK_I, Q => n_2388
                           , QN => n657);
   KEY_EXPAN0_reg_7_2_inst : FD1 port map( D => n4725, CP => CLK_I, Q => n_2389
                           , QN => n1735);
   KEY_EXPAN0_reg_6_2_inst : FD1 port map( D => n4724, CP => CLK_I, Q => n_2390
                           , QN => n664);
   KEY_EXPAN0_reg_5_2_inst : FD1 port map( D => n4723, CP => CLK_I, Q => n_2391
                           , QN => n1734);
   KEY_EXPAN0_reg_4_2_inst : FD1 port map( D => n4722, CP => CLK_I, Q => n_2392
                           , QN => n663);
   KEY_EXPAN0_reg_3_2_inst : FD1 port map( D => n4721, CP => CLK_I, Q => n_2393
                           , QN => n1733);
   KEY_EXPAN0_reg_2_2_inst : FD1 port map( D => n4720, CP => CLK_I, Q => n_2394
                           , QN => n662);
   KEY_EXPAN0_reg_1_2_inst : FD1 port map( D => n4719, CP => CLK_I, Q => n_2395
                           , QN => n1732);
   KEY_EXPAN0_reg_0_2_inst : FD1 port map( D => n4718, CP => CLK_I, Q => n_2396
                           , QN => n661);
   v_KEY_COL_OUT0_reg_2_inst : FD1 port map( D => n4560, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_2_port, QN => n1052);
   v_TEMP_VECTOR_reg_26_inst : FD1 port map( D => n6669, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_26_port, QN => n_2397);
   KEY_EXPAN0_reg_63_26_inst : FD1 port map( D => n6317, CP => CLK_I, Q => 
                           n_2398, QN => n1771);
   KEY_EXPAN0_reg_62_26_inst : FD1 port map( D => n6316, CP => CLK_I, Q => 
                           n_2399, QN => n700);
   KEY_EXPAN0_reg_61_26_inst : FD1 port map( D => n6315, CP => CLK_I, Q => 
                           n_2400, QN => n1770);
   KEY_EXPAN0_reg_60_26_inst : FD1 port map( D => n6314, CP => CLK_I, Q => 
                           n_2401, QN => n699);
   KEY_EXPAN0_reg_59_26_inst : FD1 port map( D => n6313, CP => CLK_I, Q => 
                           n_2402, QN => n1769);
   KEY_EXPAN0_reg_58_26_inst : FD1 port map( D => n6312, CP => CLK_I, Q => 
                           n_2403, QN => n698);
   KEY_EXPAN0_reg_57_26_inst : FD1 port map( D => n6311, CP => CLK_I, Q => 
                           n_2404, QN => n1768);
   KEY_EXPAN0_reg_56_26_inst : FD1 port map( D => n6310, CP => CLK_I, Q => 
                           n_2405, QN => n697);
   KEY_EXPAN0_reg_55_26_inst : FD1 port map( D => n6309, CP => CLK_I, Q => 
                           n_2406, QN => n1775);
   KEY_EXPAN0_reg_54_26_inst : FD1 port map( D => n6308, CP => CLK_I, Q => 
                           n_2407, QN => n704);
   KEY_EXPAN0_reg_53_26_inst : FD1 port map( D => n6307, CP => CLK_I, Q => 
                           n_2408, QN => n1774);
   KEY_EXPAN0_reg_52_26_inst : FD1 port map( D => n6306, CP => CLK_I, Q => 
                           n_2409, QN => n703);
   KEY_EXPAN0_reg_51_26_inst : FD1 port map( D => n6305, CP => CLK_I, Q => 
                           n_2410, QN => n1773);
   KEY_EXPAN0_reg_50_26_inst : FD1 port map( D => n6304, CP => CLK_I, Q => 
                           n_2411, QN => n702);
   KEY_EXPAN0_reg_49_26_inst : FD1 port map( D => n6303, CP => CLK_I, Q => 
                           n_2412, QN => n1772);
   KEY_EXPAN0_reg_48_26_inst : FD1 port map( D => n6302, CP => CLK_I, Q => 
                           n_2413, QN => n701);
   KEY_EXPAN0_reg_47_26_inst : FD1 port map( D => n6301, CP => CLK_I, Q => 
                           n_2414, QN => n1779);
   KEY_EXPAN0_reg_46_26_inst : FD1 port map( D => n6300, CP => CLK_I, Q => 
                           n_2415, QN => n708);
   KEY_EXPAN0_reg_45_26_inst : FD1 port map( D => n6299, CP => CLK_I, Q => 
                           n_2416, QN => n1778);
   KEY_EXPAN0_reg_44_26_inst : FD1 port map( D => n6298, CP => CLK_I, Q => 
                           n_2417, QN => n707);
   KEY_EXPAN0_reg_43_26_inst : FD1 port map( D => n6297, CP => CLK_I, Q => 
                           n_2418, QN => n1777);
   KEY_EXPAN0_reg_42_26_inst : FD1 port map( D => n6296, CP => CLK_I, Q => 
                           n_2419, QN => n706);
   KEY_EXPAN0_reg_41_26_inst : FD1 port map( D => n6295, CP => CLK_I, Q => 
                           n_2420, QN => n1776);
   KEY_EXPAN0_reg_40_26_inst : FD1 port map( D => n6294, CP => CLK_I, Q => 
                           n_2421, QN => n705);
   KEY_EXPAN0_reg_39_26_inst : FD1 port map( D => n6293, CP => CLK_I, Q => 
                           n_2422, QN => n1783);
   KEY_EXPAN0_reg_38_26_inst : FD1 port map( D => n6292, CP => CLK_I, Q => 
                           n_2423, QN => n712);
   KEY_EXPAN0_reg_37_26_inst : FD1 port map( D => n6291, CP => CLK_I, Q => 
                           n_2424, QN => n1782);
   KEY_EXPAN0_reg_36_26_inst : FD1 port map( D => n6290, CP => CLK_I, Q => 
                           n_2425, QN => n711);
   KEY_EXPAN0_reg_35_26_inst : FD1 port map( D => n6289, CP => CLK_I, Q => 
                           n_2426, QN => n1781);
   KEY_EXPAN0_reg_34_26_inst : FD1 port map( D => n6288, CP => CLK_I, Q => 
                           n_2427, QN => n710);
   KEY_EXPAN0_reg_33_26_inst : FD1 port map( D => n6287, CP => CLK_I, Q => 
                           n_2428, QN => n1780);
   KEY_EXPAN0_reg_32_26_inst : FD1 port map( D => n6286, CP => CLK_I, Q => 
                           n_2429, QN => n709);
   KEY_EXPAN0_reg_31_26_inst : FD1 port map( D => n6285, CP => CLK_I, Q => 
                           n_2430, QN => n1755);
   KEY_EXPAN0_reg_30_26_inst : FD1 port map( D => n6284, CP => CLK_I, Q => 
                           n_2431, QN => n684);
   KEY_EXPAN0_reg_29_26_inst : FD1 port map( D => n6283, CP => CLK_I, Q => 
                           n_2432, QN => n1754);
   KEY_EXPAN0_reg_28_26_inst : FD1 port map( D => n6282, CP => CLK_I, Q => 
                           n_2433, QN => n683);
   KEY_EXPAN0_reg_27_26_inst : FD1 port map( D => n6281, CP => CLK_I, Q => 
                           n_2434, QN => n1753);
   KEY_EXPAN0_reg_26_26_inst : FD1 port map( D => n6280, CP => CLK_I, Q => 
                           n_2435, QN => n682);
   KEY_EXPAN0_reg_25_26_inst : FD1 port map( D => n6279, CP => CLK_I, Q => 
                           n_2436, QN => n1752);
   KEY_EXPAN0_reg_24_26_inst : FD1 port map( D => n6278, CP => CLK_I, Q => 
                           n_2437, QN => n681);
   KEY_EXPAN0_reg_23_26_inst : FD1 port map( D => n6277, CP => CLK_I, Q => 
                           n_2438, QN => n1759);
   KEY_EXPAN0_reg_22_26_inst : FD1 port map( D => n6276, CP => CLK_I, Q => 
                           n_2439, QN => n688);
   KEY_EXPAN0_reg_21_26_inst : FD1 port map( D => n6275, CP => CLK_I, Q => 
                           n_2440, QN => n1758);
   KEY_EXPAN0_reg_20_26_inst : FD1 port map( D => n6274, CP => CLK_I, Q => 
                           n_2441, QN => n687);
   KEY_EXPAN0_reg_19_26_inst : FD1 port map( D => n6273, CP => CLK_I, Q => 
                           n_2442, QN => n1757);
   KEY_EXPAN0_reg_18_26_inst : FD1 port map( D => n6272, CP => CLK_I, Q => 
                           n_2443, QN => n686);
   KEY_EXPAN0_reg_17_26_inst : FD1 port map( D => n6271, CP => CLK_I, Q => 
                           n_2444, QN => n1756);
   KEY_EXPAN0_reg_16_26_inst : FD1 port map( D => n6270, CP => CLK_I, Q => 
                           n_2445, QN => n685);
   KEY_EXPAN0_reg_15_26_inst : FD1 port map( D => n6269, CP => CLK_I, Q => 
                           n_2446, QN => n1763);
   KEY_EXPAN0_reg_14_26_inst : FD1 port map( D => n6268, CP => CLK_I, Q => 
                           n_2447, QN => n692);
   KEY_EXPAN0_reg_13_26_inst : FD1 port map( D => n6267, CP => CLK_I, Q => 
                           n_2448, QN => n1762);
   KEY_EXPAN0_reg_12_26_inst : FD1 port map( D => n6266, CP => CLK_I, Q => 
                           n_2449, QN => n691);
   KEY_EXPAN0_reg_11_26_inst : FD1 port map( D => n6265, CP => CLK_I, Q => 
                           n_2450, QN => n1761);
   KEY_EXPAN0_reg_10_26_inst : FD1 port map( D => n6264, CP => CLK_I, Q => 
                           n_2451, QN => n690);
   KEY_EXPAN0_reg_9_26_inst : FD1 port map( D => n6263, CP => CLK_I, Q => 
                           n_2452, QN => n1760);
   KEY_EXPAN0_reg_8_26_inst : FD1 port map( D => n6262, CP => CLK_I, Q => 
                           n_2453, QN => n689);
   KEY_EXPAN0_reg_7_26_inst : FD1 port map( D => n6261, CP => CLK_I, Q => 
                           n_2454, QN => n1767);
   KEY_EXPAN0_reg_6_26_inst : FD1 port map( D => n6260, CP => CLK_I, Q => 
                           n_2455, QN => n696);
   KEY_EXPAN0_reg_5_26_inst : FD1 port map( D => n6259, CP => CLK_I, Q => 
                           n_2456, QN => n1766);
   KEY_EXPAN0_reg_4_26_inst : FD1 port map( D => n6258, CP => CLK_I, Q => 
                           n_2457, QN => n695);
   KEY_EXPAN0_reg_3_26_inst : FD1 port map( D => n6257, CP => CLK_I, Q => 
                           n_2458, QN => n1765);
   KEY_EXPAN0_reg_2_26_inst : FD1 port map( D => n6256, CP => CLK_I, Q => 
                           n_2459, QN => n694);
   KEY_EXPAN0_reg_1_26_inst : FD1 port map( D => n6255, CP => CLK_I, Q => 
                           n_2460, QN => n1764);
   KEY_EXPAN0_reg_0_26_inst : FD1 port map( D => n6254, CP => CLK_I, Q => 
                           n_2461, QN => n693);
   v_KEY_COL_OUT0_reg_26_inst : FD1 port map( D => n4559, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_26_port, QN => n1056);
   v_TEMP_VECTOR_reg_18_inst : FD1 port map( D => n6677, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_18_port, QN => n_2462);
   KEY_EXPAN0_reg_63_18_inst : FD1 port map( D => n5805, CP => CLK_I, Q => 
                           n_2463, QN => n1803);
   KEY_EXPAN0_reg_62_18_inst : FD1 port map( D => n5804, CP => CLK_I, Q => 
                           n_2464, QN => n732);
   KEY_EXPAN0_reg_61_18_inst : FD1 port map( D => n5803, CP => CLK_I, Q => 
                           n_2465, QN => n1802);
   KEY_EXPAN0_reg_60_18_inst : FD1 port map( D => n5802, CP => CLK_I, Q => 
                           n_2466, QN => n731);
   KEY_EXPAN0_reg_59_18_inst : FD1 port map( D => n5801, CP => CLK_I, Q => 
                           n_2467, QN => n1801);
   KEY_EXPAN0_reg_58_18_inst : FD1 port map( D => n5800, CP => CLK_I, Q => 
                           n_2468, QN => n730);
   KEY_EXPAN0_reg_57_18_inst : FD1 port map( D => n5799, CP => CLK_I, Q => 
                           n_2469, QN => n1800);
   KEY_EXPAN0_reg_56_18_inst : FD1 port map( D => n5798, CP => CLK_I, Q => 
                           n_2470, QN => n729);
   KEY_EXPAN0_reg_55_18_inst : FD1 port map( D => n5797, CP => CLK_I, Q => 
                           n_2471, QN => n1807);
   KEY_EXPAN0_reg_54_18_inst : FD1 port map( D => n5796, CP => CLK_I, Q => 
                           n_2472, QN => n736);
   KEY_EXPAN0_reg_53_18_inst : FD1 port map( D => n5795, CP => CLK_I, Q => 
                           n_2473, QN => n1806);
   KEY_EXPAN0_reg_52_18_inst : FD1 port map( D => n5794, CP => CLK_I, Q => 
                           n_2474, QN => n735);
   KEY_EXPAN0_reg_51_18_inst : FD1 port map( D => n5793, CP => CLK_I, Q => 
                           n_2475, QN => n1805);
   KEY_EXPAN0_reg_50_18_inst : FD1 port map( D => n5792, CP => CLK_I, Q => 
                           n_2476, QN => n734);
   KEY_EXPAN0_reg_49_18_inst : FD1 port map( D => n5791, CP => CLK_I, Q => 
                           n_2477, QN => n1804);
   KEY_EXPAN0_reg_48_18_inst : FD1 port map( D => n5790, CP => CLK_I, Q => 
                           n_2478, QN => n733);
   KEY_EXPAN0_reg_47_18_inst : FD1 port map( D => n5789, CP => CLK_I, Q => 
                           n_2479, QN => n1811);
   KEY_EXPAN0_reg_46_18_inst : FD1 port map( D => n5788, CP => CLK_I, Q => 
                           n_2480, QN => n740);
   KEY_EXPAN0_reg_45_18_inst : FD1 port map( D => n5787, CP => CLK_I, Q => 
                           n_2481, QN => n1810);
   KEY_EXPAN0_reg_44_18_inst : FD1 port map( D => n5786, CP => CLK_I, Q => 
                           n_2482, QN => n739);
   KEY_EXPAN0_reg_43_18_inst : FD1 port map( D => n5785, CP => CLK_I, Q => 
                           n_2483, QN => n1809);
   KEY_EXPAN0_reg_42_18_inst : FD1 port map( D => n5784, CP => CLK_I, Q => 
                           n_2484, QN => n738);
   KEY_EXPAN0_reg_41_18_inst : FD1 port map( D => n5783, CP => CLK_I, Q => 
                           n_2485, QN => n1808);
   KEY_EXPAN0_reg_40_18_inst : FD1 port map( D => n5782, CP => CLK_I, Q => 
                           n_2486, QN => n737);
   KEY_EXPAN0_reg_39_18_inst : FD1 port map( D => n5781, CP => CLK_I, Q => 
                           n_2487, QN => n1815);
   KEY_EXPAN0_reg_38_18_inst : FD1 port map( D => n5780, CP => CLK_I, Q => 
                           n_2488, QN => n744);
   KEY_EXPAN0_reg_37_18_inst : FD1 port map( D => n5779, CP => CLK_I, Q => 
                           n_2489, QN => n1814);
   KEY_EXPAN0_reg_36_18_inst : FD1 port map( D => n5778, CP => CLK_I, Q => 
                           n_2490, QN => n743);
   KEY_EXPAN0_reg_35_18_inst : FD1 port map( D => n5777, CP => CLK_I, Q => 
                           n_2491, QN => n1813);
   KEY_EXPAN0_reg_34_18_inst : FD1 port map( D => n5776, CP => CLK_I, Q => 
                           n_2492, QN => n742);
   KEY_EXPAN0_reg_33_18_inst : FD1 port map( D => n5775, CP => CLK_I, Q => 
                           n_2493, QN => n1812);
   KEY_EXPAN0_reg_32_18_inst : FD1 port map( D => n5774, CP => CLK_I, Q => 
                           n_2494, QN => n741);
   KEY_EXPAN0_reg_31_18_inst : FD1 port map( D => n5773, CP => CLK_I, Q => 
                           n_2495, QN => n1787);
   KEY_EXPAN0_reg_30_18_inst : FD1 port map( D => n5772, CP => CLK_I, Q => 
                           n_2496, QN => n716);
   KEY_EXPAN0_reg_29_18_inst : FD1 port map( D => n5771, CP => CLK_I, Q => 
                           n_2497, QN => n1786);
   KEY_EXPAN0_reg_28_18_inst : FD1 port map( D => n5770, CP => CLK_I, Q => 
                           n_2498, QN => n715);
   KEY_EXPAN0_reg_27_18_inst : FD1 port map( D => n5769, CP => CLK_I, Q => 
                           n_2499, QN => n1785);
   KEY_EXPAN0_reg_26_18_inst : FD1 port map( D => n5768, CP => CLK_I, Q => 
                           n_2500, QN => n714);
   KEY_EXPAN0_reg_25_18_inst : FD1 port map( D => n5767, CP => CLK_I, Q => 
                           n_2501, QN => n1784);
   KEY_EXPAN0_reg_24_18_inst : FD1 port map( D => n5766, CP => CLK_I, Q => 
                           n_2502, QN => n713);
   KEY_EXPAN0_reg_23_18_inst : FD1 port map( D => n5765, CP => CLK_I, Q => 
                           n_2503, QN => n1791);
   KEY_EXPAN0_reg_22_18_inst : FD1 port map( D => n5764, CP => CLK_I, Q => 
                           n_2504, QN => n720);
   KEY_EXPAN0_reg_21_18_inst : FD1 port map( D => n5763, CP => CLK_I, Q => 
                           n_2505, QN => n1790);
   KEY_EXPAN0_reg_20_18_inst : FD1 port map( D => n5762, CP => CLK_I, Q => 
                           n_2506, QN => n719);
   KEY_EXPAN0_reg_19_18_inst : FD1 port map( D => n5761, CP => CLK_I, Q => 
                           n_2507, QN => n1789);
   KEY_EXPAN0_reg_18_18_inst : FD1 port map( D => n5760, CP => CLK_I, Q => 
                           n_2508, QN => n718);
   KEY_EXPAN0_reg_17_18_inst : FD1 port map( D => n5759, CP => CLK_I, Q => 
                           n_2509, QN => n1788);
   KEY_EXPAN0_reg_16_18_inst : FD1 port map( D => n5758, CP => CLK_I, Q => 
                           n_2510, QN => n717);
   KEY_EXPAN0_reg_15_18_inst : FD1 port map( D => n5757, CP => CLK_I, Q => 
                           n_2511, QN => n1795);
   KEY_EXPAN0_reg_14_18_inst : FD1 port map( D => n5756, CP => CLK_I, Q => 
                           n_2512, QN => n724);
   KEY_EXPAN0_reg_13_18_inst : FD1 port map( D => n5755, CP => CLK_I, Q => 
                           n_2513, QN => n1794);
   KEY_EXPAN0_reg_12_18_inst : FD1 port map( D => n5754, CP => CLK_I, Q => 
                           n_2514, QN => n723);
   KEY_EXPAN0_reg_11_18_inst : FD1 port map( D => n5753, CP => CLK_I, Q => 
                           n_2515, QN => n1793);
   KEY_EXPAN0_reg_10_18_inst : FD1 port map( D => n5752, CP => CLK_I, Q => 
                           n_2516, QN => n722);
   KEY_EXPAN0_reg_9_18_inst : FD1 port map( D => n5751, CP => CLK_I, Q => 
                           n_2517, QN => n1792);
   KEY_EXPAN0_reg_8_18_inst : FD1 port map( D => n5750, CP => CLK_I, Q => 
                           n_2518, QN => n721);
   KEY_EXPAN0_reg_7_18_inst : FD1 port map( D => n5749, CP => CLK_I, Q => 
                           n_2519, QN => n1799);
   KEY_EXPAN0_reg_6_18_inst : FD1 port map( D => n5748, CP => CLK_I, Q => 
                           n_2520, QN => n728);
   KEY_EXPAN0_reg_5_18_inst : FD1 port map( D => n5747, CP => CLK_I, Q => 
                           n_2521, QN => n1798);
   KEY_EXPAN0_reg_4_18_inst : FD1 port map( D => n5746, CP => CLK_I, Q => 
                           n_2522, QN => n727);
   KEY_EXPAN0_reg_3_18_inst : FD1 port map( D => n5745, CP => CLK_I, Q => 
                           n_2523, QN => n1797);
   KEY_EXPAN0_reg_2_18_inst : FD1 port map( D => n5744, CP => CLK_I, Q => 
                           n_2524, QN => n726);
   KEY_EXPAN0_reg_1_18_inst : FD1 port map( D => n5743, CP => CLK_I, Q => 
                           n_2525, QN => n1796);
   KEY_EXPAN0_reg_0_18_inst : FD1 port map( D => n5742, CP => CLK_I, Q => 
                           n_2526, QN => n725);
   v_KEY_COL_OUT0_reg_18_inst : FD1 port map( D => n4558, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_18_port, QN => n1065);
   v_TEMP_VECTOR_reg_10_inst : FD1 port map( D => n6685, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_10_port, QN => n_2527);
   KEY_EXPAN0_reg_63_10_inst : FD1 port map( D => n5293, CP => CLK_I, Q => 
                           n_2528, QN => n1835);
   KEY_EXPAN0_reg_62_10_inst : FD1 port map( D => n5292, CP => CLK_I, Q => 
                           n_2529, QN => n764);
   KEY_EXPAN0_reg_61_10_inst : FD1 port map( D => n5291, CP => CLK_I, Q => 
                           n_2530, QN => n1834);
   KEY_EXPAN0_reg_60_10_inst : FD1 port map( D => n5290, CP => CLK_I, Q => 
                           n_2531, QN => n763);
   KEY_EXPAN0_reg_59_10_inst : FD1 port map( D => n5289, CP => CLK_I, Q => 
                           n_2532, QN => n1833);
   KEY_EXPAN0_reg_58_10_inst : FD1 port map( D => n5288, CP => CLK_I, Q => 
                           n_2533, QN => n762);
   KEY_EXPAN0_reg_57_10_inst : FD1 port map( D => n5287, CP => CLK_I, Q => 
                           n_2534, QN => n1832);
   KEY_EXPAN0_reg_56_10_inst : FD1 port map( D => n5286, CP => CLK_I, Q => 
                           n_2535, QN => n761);
   KEY_EXPAN0_reg_55_10_inst : FD1 port map( D => n5285, CP => CLK_I, Q => 
                           n_2536, QN => n1839);
   KEY_EXPAN0_reg_54_10_inst : FD1 port map( D => n5284, CP => CLK_I, Q => 
                           n_2537, QN => n768);
   KEY_EXPAN0_reg_53_10_inst : FD1 port map( D => n5283, CP => CLK_I, Q => 
                           n_2538, QN => n1838);
   KEY_EXPAN0_reg_52_10_inst : FD1 port map( D => n5282, CP => CLK_I, Q => 
                           n_2539, QN => n767);
   KEY_EXPAN0_reg_51_10_inst : FD1 port map( D => n5281, CP => CLK_I, Q => 
                           n_2540, QN => n1837);
   KEY_EXPAN0_reg_50_10_inst : FD1 port map( D => n5280, CP => CLK_I, Q => 
                           n_2541, QN => n766);
   KEY_EXPAN0_reg_49_10_inst : FD1 port map( D => n5279, CP => CLK_I, Q => 
                           n_2542, QN => n1836);
   KEY_EXPAN0_reg_48_10_inst : FD1 port map( D => n5278, CP => CLK_I, Q => 
                           n_2543, QN => n765);
   KEY_EXPAN0_reg_47_10_inst : FD1 port map( D => n5277, CP => CLK_I, Q => 
                           n_2544, QN => n1843);
   KEY_EXPAN0_reg_46_10_inst : FD1 port map( D => n5276, CP => CLK_I, Q => 
                           n_2545, QN => n772);
   KEY_EXPAN0_reg_45_10_inst : FD1 port map( D => n5275, CP => CLK_I, Q => 
                           n_2546, QN => n1842);
   KEY_EXPAN0_reg_44_10_inst : FD1 port map( D => n5274, CP => CLK_I, Q => 
                           n_2547, QN => n771);
   KEY_EXPAN0_reg_43_10_inst : FD1 port map( D => n5273, CP => CLK_I, Q => 
                           n_2548, QN => n1841);
   KEY_EXPAN0_reg_42_10_inst : FD1 port map( D => n5272, CP => CLK_I, Q => 
                           n_2549, QN => n770);
   KEY_EXPAN0_reg_41_10_inst : FD1 port map( D => n5271, CP => CLK_I, Q => 
                           n_2550, QN => n1840);
   KEY_EXPAN0_reg_40_10_inst : FD1 port map( D => n5270, CP => CLK_I, Q => 
                           n_2551, QN => n769);
   KEY_EXPAN0_reg_39_10_inst : FD1 port map( D => n5269, CP => CLK_I, Q => 
                           n_2552, QN => n1847);
   KEY_EXPAN0_reg_38_10_inst : FD1 port map( D => n5268, CP => CLK_I, Q => 
                           n_2553, QN => n776);
   KEY_EXPAN0_reg_37_10_inst : FD1 port map( D => n5267, CP => CLK_I, Q => 
                           n_2554, QN => n1846);
   KEY_EXPAN0_reg_36_10_inst : FD1 port map( D => n5266, CP => CLK_I, Q => 
                           n_2555, QN => n775);
   KEY_EXPAN0_reg_35_10_inst : FD1 port map( D => n5265, CP => CLK_I, Q => 
                           n_2556, QN => n1845);
   KEY_EXPAN0_reg_34_10_inst : FD1 port map( D => n5264, CP => CLK_I, Q => 
                           n_2557, QN => n774);
   KEY_EXPAN0_reg_33_10_inst : FD1 port map( D => n5263, CP => CLK_I, Q => 
                           n_2558, QN => n1844);
   KEY_EXPAN0_reg_32_10_inst : FD1 port map( D => n5262, CP => CLK_I, Q => 
                           n_2559, QN => n773);
   KEY_EXPAN0_reg_31_10_inst : FD1 port map( D => n5261, CP => CLK_I, Q => 
                           n_2560, QN => n1819);
   KEY_EXPAN0_reg_30_10_inst : FD1 port map( D => n5260, CP => CLK_I, Q => 
                           n_2561, QN => n748);
   KEY_EXPAN0_reg_29_10_inst : FD1 port map( D => n5259, CP => CLK_I, Q => 
                           n_2562, QN => n1818);
   KEY_EXPAN0_reg_28_10_inst : FD1 port map( D => n5258, CP => CLK_I, Q => 
                           n_2563, QN => n747);
   KEY_EXPAN0_reg_27_10_inst : FD1 port map( D => n5257, CP => CLK_I, Q => 
                           n_2564, QN => n1817);
   KEY_EXPAN0_reg_26_10_inst : FD1 port map( D => n5256, CP => CLK_I, Q => 
                           n_2565, QN => n746);
   KEY_EXPAN0_reg_25_10_inst : FD1 port map( D => n5255, CP => CLK_I, Q => 
                           n_2566, QN => n1816);
   KEY_EXPAN0_reg_24_10_inst : FD1 port map( D => n5254, CP => CLK_I, Q => 
                           n_2567, QN => n745);
   KEY_EXPAN0_reg_23_10_inst : FD1 port map( D => n5253, CP => CLK_I, Q => 
                           n_2568, QN => n1823);
   KEY_EXPAN0_reg_22_10_inst : FD1 port map( D => n5252, CP => CLK_I, Q => 
                           n_2569, QN => n752);
   KEY_EXPAN0_reg_21_10_inst : FD1 port map( D => n5251, CP => CLK_I, Q => 
                           n_2570, QN => n1822);
   KEY_EXPAN0_reg_20_10_inst : FD1 port map( D => n5250, CP => CLK_I, Q => 
                           n_2571, QN => n751);
   KEY_EXPAN0_reg_19_10_inst : FD1 port map( D => n5249, CP => CLK_I, Q => 
                           n_2572, QN => n1821);
   KEY_EXPAN0_reg_18_10_inst : FD1 port map( D => n5248, CP => CLK_I, Q => 
                           n_2573, QN => n750);
   KEY_EXPAN0_reg_17_10_inst : FD1 port map( D => n5247, CP => CLK_I, Q => 
                           n_2574, QN => n1820);
   KEY_EXPAN0_reg_16_10_inst : FD1 port map( D => n5246, CP => CLK_I, Q => 
                           n_2575, QN => n749);
   KEY_EXPAN0_reg_15_10_inst : FD1 port map( D => n5245, CP => CLK_I, Q => 
                           n_2576, QN => n1827);
   KEY_EXPAN0_reg_14_10_inst : FD1 port map( D => n5244, CP => CLK_I, Q => 
                           n_2577, QN => n756);
   KEY_EXPAN0_reg_13_10_inst : FD1 port map( D => n5243, CP => CLK_I, Q => 
                           n_2578, QN => n1826);
   KEY_EXPAN0_reg_12_10_inst : FD1 port map( D => n5242, CP => CLK_I, Q => 
                           n_2579, QN => n755);
   KEY_EXPAN0_reg_11_10_inst : FD1 port map( D => n5241, CP => CLK_I, Q => 
                           n_2580, QN => n1825);
   KEY_EXPAN0_reg_10_10_inst : FD1 port map( D => n5240, CP => CLK_I, Q => 
                           n_2581, QN => n754);
   KEY_EXPAN0_reg_9_10_inst : FD1 port map( D => n5239, CP => CLK_I, Q => 
                           n_2582, QN => n1824);
   KEY_EXPAN0_reg_8_10_inst : FD1 port map( D => n5238, CP => CLK_I, Q => 
                           n_2583, QN => n753);
   KEY_EXPAN0_reg_7_10_inst : FD1 port map( D => n5237, CP => CLK_I, Q => 
                           n_2584, QN => n1831);
   KEY_EXPAN0_reg_6_10_inst : FD1 port map( D => n5236, CP => CLK_I, Q => 
                           n_2585, QN => n760);
   KEY_EXPAN0_reg_5_10_inst : FD1 port map( D => n5235, CP => CLK_I, Q => 
                           n_2586, QN => n1830);
   KEY_EXPAN0_reg_4_10_inst : FD1 port map( D => n5234, CP => CLK_I, Q => 
                           n_2587, QN => n759);
   KEY_EXPAN0_reg_3_10_inst : FD1 port map( D => n5233, CP => CLK_I, Q => 
                           n_2588, QN => n1829);
   KEY_EXPAN0_reg_2_10_inst : FD1 port map( D => n5232, CP => CLK_I, Q => 
                           n_2589, QN => n758);
   KEY_EXPAN0_reg_1_10_inst : FD1 port map( D => n5231, CP => CLK_I, Q => 
                           n_2590, QN => n1828);
   KEY_EXPAN0_reg_0_10_inst : FD1 port map( D => n5230, CP => CLK_I, Q => 
                           n_2591, QN => n757);
   v_KEY_COL_OUT0_reg_10_inst : FD1 port map( D => n4557, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_10_port, QN => n1073);
   v_TEMP_VECTOR_reg_1_inst : FD1 port map( D => n6694, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_1_port, QN => n_2592);
   KEY_EXPAN0_reg_63_1_inst : FD1 port map( D => n4717, CP => CLK_I, Q => 
                           n_2593, QN => n1867);
   KEY_EXPAN0_reg_62_1_inst : FD1 port map( D => n4716, CP => CLK_I, Q => 
                           n_2594, QN => n796);
   KEY_EXPAN0_reg_61_1_inst : FD1 port map( D => n4715, CP => CLK_I, Q => 
                           n_2595, QN => n1866);
   KEY_EXPAN0_reg_60_1_inst : FD1 port map( D => n4714, CP => CLK_I, Q => 
                           n_2596, QN => n795);
   KEY_EXPAN0_reg_59_1_inst : FD1 port map( D => n4713, CP => CLK_I, Q => 
                           n_2597, QN => n1865);
   KEY_EXPAN0_reg_58_1_inst : FD1 port map( D => n4712, CP => CLK_I, Q => 
                           n_2598, QN => n794);
   KEY_EXPAN0_reg_57_1_inst : FD1 port map( D => n4711, CP => CLK_I, Q => 
                           n_2599, QN => n1864);
   KEY_EXPAN0_reg_56_1_inst : FD1 port map( D => n4710, CP => CLK_I, Q => 
                           n_2600, QN => n793);
   KEY_EXPAN0_reg_55_1_inst : FD1 port map( D => n4709, CP => CLK_I, Q => 
                           n_2601, QN => n1871);
   KEY_EXPAN0_reg_54_1_inst : FD1 port map( D => n4708, CP => CLK_I, Q => 
                           n_2602, QN => n800);
   KEY_EXPAN0_reg_53_1_inst : FD1 port map( D => n4707, CP => CLK_I, Q => 
                           n_2603, QN => n1870);
   KEY_EXPAN0_reg_52_1_inst : FD1 port map( D => n4706, CP => CLK_I, Q => 
                           n_2604, QN => n799);
   KEY_EXPAN0_reg_51_1_inst : FD1 port map( D => n4705, CP => CLK_I, Q => 
                           n_2605, QN => n1869);
   KEY_EXPAN0_reg_50_1_inst : FD1 port map( D => n4704, CP => CLK_I, Q => 
                           n_2606, QN => n798);
   KEY_EXPAN0_reg_49_1_inst : FD1 port map( D => n4703, CP => CLK_I, Q => 
                           n_2607, QN => n1868);
   KEY_EXPAN0_reg_48_1_inst : FD1 port map( D => n4702, CP => CLK_I, Q => 
                           n_2608, QN => n797);
   KEY_EXPAN0_reg_47_1_inst : FD1 port map( D => n4701, CP => CLK_I, Q => 
                           n_2609, QN => n1875);
   KEY_EXPAN0_reg_46_1_inst : FD1 port map( D => n4700, CP => CLK_I, Q => 
                           n_2610, QN => n804);
   KEY_EXPAN0_reg_45_1_inst : FD1 port map( D => n4699, CP => CLK_I, Q => 
                           n_2611, QN => n1874);
   KEY_EXPAN0_reg_44_1_inst : FD1 port map( D => n4698, CP => CLK_I, Q => 
                           n_2612, QN => n803);
   KEY_EXPAN0_reg_43_1_inst : FD1 port map( D => n4697, CP => CLK_I, Q => 
                           n_2613, QN => n1873);
   KEY_EXPAN0_reg_42_1_inst : FD1 port map( D => n4696, CP => CLK_I, Q => 
                           n_2614, QN => n802);
   KEY_EXPAN0_reg_41_1_inst : FD1 port map( D => n4695, CP => CLK_I, Q => 
                           n_2615, QN => n1872);
   KEY_EXPAN0_reg_40_1_inst : FD1 port map( D => n4694, CP => CLK_I, Q => 
                           n_2616, QN => n801);
   KEY_EXPAN0_reg_39_1_inst : FD1 port map( D => n4693, CP => CLK_I, Q => 
                           n_2617, QN => n1879);
   KEY_EXPAN0_reg_38_1_inst : FD1 port map( D => n4692, CP => CLK_I, Q => 
                           n_2618, QN => n808);
   KEY_EXPAN0_reg_37_1_inst : FD1 port map( D => n4691, CP => CLK_I, Q => 
                           n_2619, QN => n1878);
   KEY_EXPAN0_reg_36_1_inst : FD1 port map( D => n4690, CP => CLK_I, Q => 
                           n_2620, QN => n807);
   KEY_EXPAN0_reg_35_1_inst : FD1 port map( D => n4689, CP => CLK_I, Q => 
                           n_2621, QN => n1877);
   KEY_EXPAN0_reg_34_1_inst : FD1 port map( D => n4688, CP => CLK_I, Q => 
                           n_2622, QN => n806);
   KEY_EXPAN0_reg_33_1_inst : FD1 port map( D => n4687, CP => CLK_I, Q => 
                           n_2623, QN => n1876);
   KEY_EXPAN0_reg_32_1_inst : FD1 port map( D => n4686, CP => CLK_I, Q => 
                           n_2624, QN => n805);
   KEY_EXPAN0_reg_31_1_inst : FD1 port map( D => n4685, CP => CLK_I, Q => 
                           n_2625, QN => n1851);
   KEY_EXPAN0_reg_30_1_inst : FD1 port map( D => n4684, CP => CLK_I, Q => 
                           n_2626, QN => n780);
   KEY_EXPAN0_reg_29_1_inst : FD1 port map( D => n4683, CP => CLK_I, Q => 
                           n_2627, QN => n1850);
   KEY_EXPAN0_reg_28_1_inst : FD1 port map( D => n4682, CP => CLK_I, Q => 
                           n_2628, QN => n779);
   KEY_EXPAN0_reg_27_1_inst : FD1 port map( D => n4681, CP => CLK_I, Q => 
                           n_2629, QN => n1849);
   KEY_EXPAN0_reg_26_1_inst : FD1 port map( D => n4680, CP => CLK_I, Q => 
                           n_2630, QN => n778);
   KEY_EXPAN0_reg_25_1_inst : FD1 port map( D => n4679, CP => CLK_I, Q => 
                           n_2631, QN => n1848);
   KEY_EXPAN0_reg_24_1_inst : FD1 port map( D => n4678, CP => CLK_I, Q => 
                           n_2632, QN => n777);
   KEY_EXPAN0_reg_23_1_inst : FD1 port map( D => n4677, CP => CLK_I, Q => 
                           n_2633, QN => n1855);
   KEY_EXPAN0_reg_22_1_inst : FD1 port map( D => n4676, CP => CLK_I, Q => 
                           n_2634, QN => n784);
   KEY_EXPAN0_reg_21_1_inst : FD1 port map( D => n4675, CP => CLK_I, Q => 
                           n_2635, QN => n1854);
   KEY_EXPAN0_reg_20_1_inst : FD1 port map( D => n4674, CP => CLK_I, Q => 
                           n_2636, QN => n783);
   KEY_EXPAN0_reg_19_1_inst : FD1 port map( D => n4673, CP => CLK_I, Q => 
                           n_2637, QN => n1853);
   KEY_EXPAN0_reg_18_1_inst : FD1 port map( D => n4672, CP => CLK_I, Q => 
                           n_2638, QN => n782);
   KEY_EXPAN0_reg_17_1_inst : FD1 port map( D => n4671, CP => CLK_I, Q => 
                           n_2639, QN => n1852);
   KEY_EXPAN0_reg_16_1_inst : FD1 port map( D => n4670, CP => CLK_I, Q => 
                           n_2640, QN => n781);
   KEY_EXPAN0_reg_15_1_inst : FD1 port map( D => n4669, CP => CLK_I, Q => 
                           n_2641, QN => n1859);
   KEY_EXPAN0_reg_14_1_inst : FD1 port map( D => n4668, CP => CLK_I, Q => 
                           n_2642, QN => n788);
   KEY_EXPAN0_reg_13_1_inst : FD1 port map( D => n4667, CP => CLK_I, Q => 
                           n_2643, QN => n1858);
   KEY_EXPAN0_reg_12_1_inst : FD1 port map( D => n4666, CP => CLK_I, Q => 
                           n_2644, QN => n787);
   KEY_EXPAN0_reg_11_1_inst : FD1 port map( D => n4665, CP => CLK_I, Q => 
                           n_2645, QN => n1857);
   KEY_EXPAN0_reg_10_1_inst : FD1 port map( D => n4664, CP => CLK_I, Q => 
                           n_2646, QN => n786);
   KEY_EXPAN0_reg_9_1_inst : FD1 port map( D => n4663, CP => CLK_I, Q => n_2647
                           , QN => n1856);
   KEY_EXPAN0_reg_8_1_inst : FD1 port map( D => n4662, CP => CLK_I, Q => n_2648
                           , QN => n785);
   KEY_EXPAN0_reg_7_1_inst : FD1 port map( D => n4661, CP => CLK_I, Q => n_2649
                           , QN => n1863);
   KEY_EXPAN0_reg_6_1_inst : FD1 port map( D => n4660, CP => CLK_I, Q => n_2650
                           , QN => n792);
   KEY_EXPAN0_reg_5_1_inst : FD1 port map( D => n4659, CP => CLK_I, Q => n_2651
                           , QN => n1862);
   KEY_EXPAN0_reg_4_1_inst : FD1 port map( D => n4658, CP => CLK_I, Q => n_2652
                           , QN => n791);
   KEY_EXPAN0_reg_3_1_inst : FD1 port map( D => n4657, CP => CLK_I, Q => n_2653
                           , QN => n1861);
   KEY_EXPAN0_reg_2_1_inst : FD1 port map( D => n4656, CP => CLK_I, Q => n_2654
                           , QN => n790);
   KEY_EXPAN0_reg_1_1_inst : FD1 port map( D => n4655, CP => CLK_I, Q => n_2655
                           , QN => n1860);
   KEY_EXPAN0_reg_0_1_inst : FD1 port map( D => n4654, CP => CLK_I, Q => n_2656
                           , QN => n789);
   v_KEY_COL_OUT0_reg_1_inst : FD1 port map( D => n4556, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_1_port, QN => n1063);
   v_TEMP_VECTOR_reg_25_inst : FD1 port map( D => n6670, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_25_port, QN => n_2657);
   KEY_EXPAN0_reg_63_25_inst : FD1 port map( D => n6253, CP => CLK_I, Q => 
                           n_2658, QN => n1899);
   KEY_EXPAN0_reg_62_25_inst : FD1 port map( D => n6252, CP => CLK_I, Q => 
                           n_2659, QN => n828);
   KEY_EXPAN0_reg_61_25_inst : FD1 port map( D => n6251, CP => CLK_I, Q => 
                           n_2660, QN => n1898);
   KEY_EXPAN0_reg_60_25_inst : FD1 port map( D => n6250, CP => CLK_I, Q => 
                           n_2661, QN => n827);
   KEY_EXPAN0_reg_59_25_inst : FD1 port map( D => n6249, CP => CLK_I, Q => 
                           n_2662, QN => n1897);
   KEY_EXPAN0_reg_58_25_inst : FD1 port map( D => n6248, CP => CLK_I, Q => 
                           n_2663, QN => n826);
   KEY_EXPAN0_reg_57_25_inst : FD1 port map( D => n6247, CP => CLK_I, Q => 
                           n_2664, QN => n1896);
   KEY_EXPAN0_reg_56_25_inst : FD1 port map( D => n6246, CP => CLK_I, Q => 
                           n_2665, QN => n825);
   KEY_EXPAN0_reg_55_25_inst : FD1 port map( D => n6245, CP => CLK_I, Q => 
                           n_2666, QN => n1903);
   KEY_EXPAN0_reg_54_25_inst : FD1 port map( D => n6244, CP => CLK_I, Q => 
                           n_2667, QN => n832);
   KEY_EXPAN0_reg_53_25_inst : FD1 port map( D => n6243, CP => CLK_I, Q => 
                           n_2668, QN => n1902);
   KEY_EXPAN0_reg_52_25_inst : FD1 port map( D => n6242, CP => CLK_I, Q => 
                           n_2669, QN => n831);
   KEY_EXPAN0_reg_51_25_inst : FD1 port map( D => n6241, CP => CLK_I, Q => 
                           n_2670, QN => n1901);
   KEY_EXPAN0_reg_50_25_inst : FD1 port map( D => n6240, CP => CLK_I, Q => 
                           n_2671, QN => n830);
   KEY_EXPAN0_reg_49_25_inst : FD1 port map( D => n6239, CP => CLK_I, Q => 
                           n_2672, QN => n1900);
   KEY_EXPAN0_reg_48_25_inst : FD1 port map( D => n6238, CP => CLK_I, Q => 
                           n_2673, QN => n829);
   KEY_EXPAN0_reg_47_25_inst : FD1 port map( D => n6237, CP => CLK_I, Q => 
                           n_2674, QN => n1907);
   KEY_EXPAN0_reg_46_25_inst : FD1 port map( D => n6236, CP => CLK_I, Q => 
                           n_2675, QN => n836);
   KEY_EXPAN0_reg_45_25_inst : FD1 port map( D => n6235, CP => CLK_I, Q => 
                           n_2676, QN => n1906);
   KEY_EXPAN0_reg_44_25_inst : FD1 port map( D => n6234, CP => CLK_I, Q => 
                           n_2677, QN => n835);
   KEY_EXPAN0_reg_43_25_inst : FD1 port map( D => n6233, CP => CLK_I, Q => 
                           n_2678, QN => n1905);
   KEY_EXPAN0_reg_42_25_inst : FD1 port map( D => n6232, CP => CLK_I, Q => 
                           n_2679, QN => n834);
   KEY_EXPAN0_reg_41_25_inst : FD1 port map( D => n6231, CP => CLK_I, Q => 
                           n_2680, QN => n1904);
   KEY_EXPAN0_reg_40_25_inst : FD1 port map( D => n6230, CP => CLK_I, Q => 
                           n_2681, QN => n833);
   KEY_EXPAN0_reg_39_25_inst : FD1 port map( D => n6229, CP => CLK_I, Q => 
                           n_2682, QN => n1911);
   KEY_EXPAN0_reg_38_25_inst : FD1 port map( D => n6228, CP => CLK_I, Q => 
                           n_2683, QN => n840);
   KEY_EXPAN0_reg_37_25_inst : FD1 port map( D => n6227, CP => CLK_I, Q => 
                           n_2684, QN => n1910);
   KEY_EXPAN0_reg_36_25_inst : FD1 port map( D => n6226, CP => CLK_I, Q => 
                           n_2685, QN => n839);
   KEY_EXPAN0_reg_35_25_inst : FD1 port map( D => n6225, CP => CLK_I, Q => 
                           n_2686, QN => n1909);
   KEY_EXPAN0_reg_34_25_inst : FD1 port map( D => n6224, CP => CLK_I, Q => 
                           n_2687, QN => n838);
   KEY_EXPAN0_reg_33_25_inst : FD1 port map( D => n6223, CP => CLK_I, Q => 
                           n_2688, QN => n1908);
   KEY_EXPAN0_reg_32_25_inst : FD1 port map( D => n6222, CP => CLK_I, Q => 
                           n_2689, QN => n837);
   KEY_EXPAN0_reg_31_25_inst : FD1 port map( D => n6221, CP => CLK_I, Q => 
                           n_2690, QN => n1883);
   KEY_EXPAN0_reg_30_25_inst : FD1 port map( D => n6220, CP => CLK_I, Q => 
                           n_2691, QN => n812);
   KEY_EXPAN0_reg_29_25_inst : FD1 port map( D => n6219, CP => CLK_I, Q => 
                           n_2692, QN => n1882);
   KEY_EXPAN0_reg_28_25_inst : FD1 port map( D => n6218, CP => CLK_I, Q => 
                           n_2693, QN => n811);
   KEY_EXPAN0_reg_27_25_inst : FD1 port map( D => n6217, CP => CLK_I, Q => 
                           n_2694, QN => n1881);
   KEY_EXPAN0_reg_26_25_inst : FD1 port map( D => n6216, CP => CLK_I, Q => 
                           n_2695, QN => n810);
   KEY_EXPAN0_reg_25_25_inst : FD1 port map( D => n6215, CP => CLK_I, Q => 
                           n_2696, QN => n1880);
   KEY_EXPAN0_reg_24_25_inst : FD1 port map( D => n6214, CP => CLK_I, Q => 
                           n_2697, QN => n809);
   KEY_EXPAN0_reg_23_25_inst : FD1 port map( D => n6213, CP => CLK_I, Q => 
                           n_2698, QN => n1887);
   KEY_EXPAN0_reg_22_25_inst : FD1 port map( D => n6212, CP => CLK_I, Q => 
                           n_2699, QN => n816);
   KEY_EXPAN0_reg_21_25_inst : FD1 port map( D => n6211, CP => CLK_I, Q => 
                           n_2700, QN => n1886);
   KEY_EXPAN0_reg_20_25_inst : FD1 port map( D => n6210, CP => CLK_I, Q => 
                           n_2701, QN => n815);
   KEY_EXPAN0_reg_19_25_inst : FD1 port map( D => n6209, CP => CLK_I, Q => 
                           n_2702, QN => n1885);
   KEY_EXPAN0_reg_18_25_inst : FD1 port map( D => n6208, CP => CLK_I, Q => 
                           n_2703, QN => n814);
   KEY_EXPAN0_reg_17_25_inst : FD1 port map( D => n6207, CP => CLK_I, Q => 
                           n_2704, QN => n1884);
   KEY_EXPAN0_reg_16_25_inst : FD1 port map( D => n6206, CP => CLK_I, Q => 
                           n_2705, QN => n813);
   KEY_EXPAN0_reg_15_25_inst : FD1 port map( D => n6205, CP => CLK_I, Q => 
                           n_2706, QN => n1891);
   KEY_EXPAN0_reg_14_25_inst : FD1 port map( D => n6204, CP => CLK_I, Q => 
                           n_2707, QN => n820);
   KEY_EXPAN0_reg_13_25_inst : FD1 port map( D => n6203, CP => CLK_I, Q => 
                           n_2708, QN => n1890);
   KEY_EXPAN0_reg_12_25_inst : FD1 port map( D => n6202, CP => CLK_I, Q => 
                           n_2709, QN => n819);
   KEY_EXPAN0_reg_11_25_inst : FD1 port map( D => n6201, CP => CLK_I, Q => 
                           n_2710, QN => n1889);
   KEY_EXPAN0_reg_10_25_inst : FD1 port map( D => n6200, CP => CLK_I, Q => 
                           n_2711, QN => n818);
   KEY_EXPAN0_reg_9_25_inst : FD1 port map( D => n6199, CP => CLK_I, Q => 
                           n_2712, QN => n1888);
   KEY_EXPAN0_reg_8_25_inst : FD1 port map( D => n6198, CP => CLK_I, Q => 
                           n_2713, QN => n817);
   KEY_EXPAN0_reg_7_25_inst : FD1 port map( D => n6197, CP => CLK_I, Q => 
                           n_2714, QN => n1895);
   KEY_EXPAN0_reg_6_25_inst : FD1 port map( D => n6196, CP => CLK_I, Q => 
                           n_2715, QN => n824);
   KEY_EXPAN0_reg_5_25_inst : FD1 port map( D => n6195, CP => CLK_I, Q => 
                           n_2716, QN => n1894);
   KEY_EXPAN0_reg_4_25_inst : FD1 port map( D => n6194, CP => CLK_I, Q => 
                           n_2717, QN => n823);
   KEY_EXPAN0_reg_3_25_inst : FD1 port map( D => n6193, CP => CLK_I, Q => 
                           n_2718, QN => n1893);
   KEY_EXPAN0_reg_2_25_inst : FD1 port map( D => n6192, CP => CLK_I, Q => 
                           n_2719, QN => n822);
   KEY_EXPAN0_reg_1_25_inst : FD1 port map( D => n6191, CP => CLK_I, Q => 
                           n_2720, QN => n1892);
   KEY_EXPAN0_reg_0_25_inst : FD1 port map( D => n6190, CP => CLK_I, Q => 
                           n_2721, QN => n821);
   v_KEY_COL_OUT0_reg_25_inst : FD1 port map( D => n4555, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_25_port, QN => n1057);
   v_TEMP_VECTOR_reg_17_inst : FD1 port map( D => n6678, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_17_port, QN => n_2722);
   KEY_EXPAN0_reg_63_17_inst : FD1 port map( D => n5741, CP => CLK_I, Q => 
                           n_2723, QN => n1931);
   KEY_EXPAN0_reg_62_17_inst : FD1 port map( D => n5740, CP => CLK_I, Q => 
                           n_2724, QN => n860);
   KEY_EXPAN0_reg_61_17_inst : FD1 port map( D => n5739, CP => CLK_I, Q => 
                           n_2725, QN => n1930);
   KEY_EXPAN0_reg_60_17_inst : FD1 port map( D => n5738, CP => CLK_I, Q => 
                           n_2726, QN => n859);
   KEY_EXPAN0_reg_59_17_inst : FD1 port map( D => n5737, CP => CLK_I, Q => 
                           n_2727, QN => n1929);
   KEY_EXPAN0_reg_58_17_inst : FD1 port map( D => n5736, CP => CLK_I, Q => 
                           n_2728, QN => n858);
   KEY_EXPAN0_reg_57_17_inst : FD1 port map( D => n5735, CP => CLK_I, Q => 
                           n_2729, QN => n1928);
   KEY_EXPAN0_reg_56_17_inst : FD1 port map( D => n5734, CP => CLK_I, Q => 
                           n_2730, QN => n857);
   KEY_EXPAN0_reg_55_17_inst : FD1 port map( D => n5733, CP => CLK_I, Q => 
                           n_2731, QN => n1935);
   KEY_EXPAN0_reg_54_17_inst : FD1 port map( D => n5732, CP => CLK_I, Q => 
                           n_2732, QN => n864);
   KEY_EXPAN0_reg_53_17_inst : FD1 port map( D => n5731, CP => CLK_I, Q => 
                           n_2733, QN => n1934);
   KEY_EXPAN0_reg_52_17_inst : FD1 port map( D => n5730, CP => CLK_I, Q => 
                           n_2734, QN => n863);
   KEY_EXPAN0_reg_51_17_inst : FD1 port map( D => n5729, CP => CLK_I, Q => 
                           n_2735, QN => n1933);
   KEY_EXPAN0_reg_50_17_inst : FD1 port map( D => n5728, CP => CLK_I, Q => 
                           n_2736, QN => n862);
   KEY_EXPAN0_reg_49_17_inst : FD1 port map( D => n5727, CP => CLK_I, Q => 
                           n_2737, QN => n1932);
   KEY_EXPAN0_reg_48_17_inst : FD1 port map( D => n5726, CP => CLK_I, Q => 
                           n_2738, QN => n861);
   KEY_EXPAN0_reg_47_17_inst : FD1 port map( D => n5725, CP => CLK_I, Q => 
                           n_2739, QN => n1939);
   KEY_EXPAN0_reg_46_17_inst : FD1 port map( D => n5724, CP => CLK_I, Q => 
                           n_2740, QN => n868);
   KEY_EXPAN0_reg_45_17_inst : FD1 port map( D => n5723, CP => CLK_I, Q => 
                           n_2741, QN => n1938);
   KEY_EXPAN0_reg_44_17_inst : FD1 port map( D => n5722, CP => CLK_I, Q => 
                           n_2742, QN => n867);
   KEY_EXPAN0_reg_43_17_inst : FD1 port map( D => n5721, CP => CLK_I, Q => 
                           n_2743, QN => n1937);
   KEY_EXPAN0_reg_42_17_inst : FD1 port map( D => n5720, CP => CLK_I, Q => 
                           n_2744, QN => n866);
   KEY_EXPAN0_reg_41_17_inst : FD1 port map( D => n5719, CP => CLK_I, Q => 
                           n_2745, QN => n1936);
   KEY_EXPAN0_reg_40_17_inst : FD1 port map( D => n5718, CP => CLK_I, Q => 
                           n_2746, QN => n865);
   KEY_EXPAN0_reg_39_17_inst : FD1 port map( D => n5717, CP => CLK_I, Q => 
                           n_2747, QN => n1943);
   KEY_EXPAN0_reg_38_17_inst : FD1 port map( D => n5716, CP => CLK_I, Q => 
                           n_2748, QN => n872);
   KEY_EXPAN0_reg_37_17_inst : FD1 port map( D => n5715, CP => CLK_I, Q => 
                           n_2749, QN => n1942);
   KEY_EXPAN0_reg_36_17_inst : FD1 port map( D => n5714, CP => CLK_I, Q => 
                           n_2750, QN => n871);
   KEY_EXPAN0_reg_35_17_inst : FD1 port map( D => n5713, CP => CLK_I, Q => 
                           n_2751, QN => n1941);
   KEY_EXPAN0_reg_34_17_inst : FD1 port map( D => n5712, CP => CLK_I, Q => 
                           n_2752, QN => n870);
   KEY_EXPAN0_reg_33_17_inst : FD1 port map( D => n5711, CP => CLK_I, Q => 
                           n_2753, QN => n1940);
   KEY_EXPAN0_reg_32_17_inst : FD1 port map( D => n5710, CP => CLK_I, Q => 
                           n_2754, QN => n869);
   KEY_EXPAN0_reg_31_17_inst : FD1 port map( D => n5709, CP => CLK_I, Q => 
                           n_2755, QN => n1915);
   KEY_EXPAN0_reg_30_17_inst : FD1 port map( D => n5708, CP => CLK_I, Q => 
                           n_2756, QN => n844);
   KEY_EXPAN0_reg_29_17_inst : FD1 port map( D => n5707, CP => CLK_I, Q => 
                           n_2757, QN => n1914);
   KEY_EXPAN0_reg_28_17_inst : FD1 port map( D => n5706, CP => CLK_I, Q => 
                           n_2758, QN => n843);
   KEY_EXPAN0_reg_27_17_inst : FD1 port map( D => n5705, CP => CLK_I, Q => 
                           n_2759, QN => n1913);
   KEY_EXPAN0_reg_26_17_inst : FD1 port map( D => n5704, CP => CLK_I, Q => 
                           n_2760, QN => n842);
   KEY_EXPAN0_reg_25_17_inst : FD1 port map( D => n5703, CP => CLK_I, Q => 
                           n_2761, QN => n1912);
   KEY_EXPAN0_reg_24_17_inst : FD1 port map( D => n5702, CP => CLK_I, Q => 
                           n_2762, QN => n841);
   KEY_EXPAN0_reg_23_17_inst : FD1 port map( D => n5701, CP => CLK_I, Q => 
                           n_2763, QN => n1919);
   KEY_EXPAN0_reg_22_17_inst : FD1 port map( D => n5700, CP => CLK_I, Q => 
                           n_2764, QN => n848);
   KEY_EXPAN0_reg_21_17_inst : FD1 port map( D => n5699, CP => CLK_I, Q => 
                           n_2765, QN => n1918);
   KEY_EXPAN0_reg_20_17_inst : FD1 port map( D => n5698, CP => CLK_I, Q => 
                           n_2766, QN => n847);
   KEY_EXPAN0_reg_19_17_inst : FD1 port map( D => n5697, CP => CLK_I, Q => 
                           n_2767, QN => n1917);
   KEY_EXPAN0_reg_18_17_inst : FD1 port map( D => n5696, CP => CLK_I, Q => 
                           n_2768, QN => n846);
   KEY_EXPAN0_reg_17_17_inst : FD1 port map( D => n5695, CP => CLK_I, Q => 
                           n_2769, QN => n1916);
   KEY_EXPAN0_reg_16_17_inst : FD1 port map( D => n5694, CP => CLK_I, Q => 
                           n_2770, QN => n845);
   KEY_EXPAN0_reg_15_17_inst : FD1 port map( D => n5693, CP => CLK_I, Q => 
                           n_2771, QN => n1923);
   KEY_EXPAN0_reg_14_17_inst : FD1 port map( D => n5692, CP => CLK_I, Q => 
                           n_2772, QN => n852);
   KEY_EXPAN0_reg_13_17_inst : FD1 port map( D => n5691, CP => CLK_I, Q => 
                           n_2773, QN => n1922);
   KEY_EXPAN0_reg_12_17_inst : FD1 port map( D => n5690, CP => CLK_I, Q => 
                           n_2774, QN => n851);
   KEY_EXPAN0_reg_11_17_inst : FD1 port map( D => n5689, CP => CLK_I, Q => 
                           n_2775, QN => n1921);
   KEY_EXPAN0_reg_10_17_inst : FD1 port map( D => n5688, CP => CLK_I, Q => 
                           n_2776, QN => n850);
   KEY_EXPAN0_reg_9_17_inst : FD1 port map( D => n5687, CP => CLK_I, Q => 
                           n_2777, QN => n1920);
   KEY_EXPAN0_reg_8_17_inst : FD1 port map( D => n5686, CP => CLK_I, Q => 
                           n_2778, QN => n849);
   KEY_EXPAN0_reg_7_17_inst : FD1 port map( D => n5685, CP => CLK_I, Q => 
                           n_2779, QN => n1927);
   KEY_EXPAN0_reg_6_17_inst : FD1 port map( D => n5684, CP => CLK_I, Q => 
                           n_2780, QN => n856);
   KEY_EXPAN0_reg_5_17_inst : FD1 port map( D => n5683, CP => CLK_I, Q => 
                           n_2781, QN => n1926);
   KEY_EXPAN0_reg_4_17_inst : FD1 port map( D => n5682, CP => CLK_I, Q => 
                           n_2782, QN => n855);
   KEY_EXPAN0_reg_3_17_inst : FD1 port map( D => n5681, CP => CLK_I, Q => 
                           n_2783, QN => n1925);
   KEY_EXPAN0_reg_2_17_inst : FD1 port map( D => n5680, CP => CLK_I, Q => 
                           n_2784, QN => n854);
   KEY_EXPAN0_reg_1_17_inst : FD1 port map( D => n5679, CP => CLK_I, Q => 
                           n_2785, QN => n1924);
   KEY_EXPAN0_reg_0_17_inst : FD1 port map( D => n5678, CP => CLK_I, Q => 
                           n_2786, QN => n853);
   v_KEY_COL_OUT0_reg_17_inst : FD1 port map( D => n4554, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_17_port, QN => n1066);
   v_TEMP_VECTOR_reg_9_inst : FD1 port map( D => n6686, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_9_port, QN => n_2787);
   KEY_EXPAN0_reg_63_9_inst : FD1 port map( D => n5229, CP => CLK_I, Q => 
                           n_2788, QN => n1963);
   KEY_EXPAN0_reg_62_9_inst : FD1 port map( D => n5228, CP => CLK_I, Q => 
                           n_2789, QN => n892);
   KEY_EXPAN0_reg_61_9_inst : FD1 port map( D => n5227, CP => CLK_I, Q => 
                           n_2790, QN => n1962);
   KEY_EXPAN0_reg_60_9_inst : FD1 port map( D => n5226, CP => CLK_I, Q => 
                           n_2791, QN => n891);
   KEY_EXPAN0_reg_59_9_inst : FD1 port map( D => n5225, CP => CLK_I, Q => 
                           n_2792, QN => n1961);
   KEY_EXPAN0_reg_58_9_inst : FD1 port map( D => n5224, CP => CLK_I, Q => 
                           n_2793, QN => n890);
   KEY_EXPAN0_reg_57_9_inst : FD1 port map( D => n5223, CP => CLK_I, Q => 
                           n_2794, QN => n1960);
   KEY_EXPAN0_reg_56_9_inst : FD1 port map( D => n5222, CP => CLK_I, Q => 
                           n_2795, QN => n889);
   KEY_EXPAN0_reg_55_9_inst : FD1 port map( D => n5221, CP => CLK_I, Q => 
                           n_2796, QN => n1967);
   KEY_EXPAN0_reg_54_9_inst : FD1 port map( D => n5220, CP => CLK_I, Q => 
                           n_2797, QN => n896);
   KEY_EXPAN0_reg_53_9_inst : FD1 port map( D => n5219, CP => CLK_I, Q => 
                           n_2798, QN => n1966);
   KEY_EXPAN0_reg_52_9_inst : FD1 port map( D => n5218, CP => CLK_I, Q => 
                           n_2799, QN => n895);
   KEY_EXPAN0_reg_51_9_inst : FD1 port map( D => n5217, CP => CLK_I, Q => 
                           n_2800, QN => n1965);
   KEY_EXPAN0_reg_50_9_inst : FD1 port map( D => n5216, CP => CLK_I, Q => 
                           n_2801, QN => n894);
   KEY_EXPAN0_reg_49_9_inst : FD1 port map( D => n5215, CP => CLK_I, Q => 
                           n_2802, QN => n1964);
   KEY_EXPAN0_reg_48_9_inst : FD1 port map( D => n5214, CP => CLK_I, Q => 
                           n_2803, QN => n893);
   KEY_EXPAN0_reg_47_9_inst : FD1 port map( D => n5213, CP => CLK_I, Q => 
                           n_2804, QN => n1971);
   KEY_EXPAN0_reg_46_9_inst : FD1 port map( D => n5212, CP => CLK_I, Q => 
                           n_2805, QN => n900);
   KEY_EXPAN0_reg_45_9_inst : FD1 port map( D => n5211, CP => CLK_I, Q => 
                           n_2806, QN => n1970);
   KEY_EXPAN0_reg_44_9_inst : FD1 port map( D => n5210, CP => CLK_I, Q => 
                           n_2807, QN => n899);
   KEY_EXPAN0_reg_43_9_inst : FD1 port map( D => n5209, CP => CLK_I, Q => 
                           n_2808, QN => n1969);
   KEY_EXPAN0_reg_42_9_inst : FD1 port map( D => n5208, CP => CLK_I, Q => 
                           n_2809, QN => n898);
   KEY_EXPAN0_reg_41_9_inst : FD1 port map( D => n5207, CP => CLK_I, Q => 
                           n_2810, QN => n1968);
   KEY_EXPAN0_reg_40_9_inst : FD1 port map( D => n5206, CP => CLK_I, Q => 
                           n_2811, QN => n897);
   KEY_EXPAN0_reg_39_9_inst : FD1 port map( D => n5205, CP => CLK_I, Q => 
                           n_2812, QN => n1975);
   KEY_EXPAN0_reg_38_9_inst : FD1 port map( D => n5204, CP => CLK_I, Q => 
                           n_2813, QN => n904);
   KEY_EXPAN0_reg_37_9_inst : FD1 port map( D => n5203, CP => CLK_I, Q => 
                           n_2814, QN => n1974);
   KEY_EXPAN0_reg_36_9_inst : FD1 port map( D => n5202, CP => CLK_I, Q => 
                           n_2815, QN => n903);
   KEY_EXPAN0_reg_35_9_inst : FD1 port map( D => n5201, CP => CLK_I, Q => 
                           n_2816, QN => n1973);
   KEY_EXPAN0_reg_34_9_inst : FD1 port map( D => n5200, CP => CLK_I, Q => 
                           n_2817, QN => n902);
   KEY_EXPAN0_reg_33_9_inst : FD1 port map( D => n5199, CP => CLK_I, Q => 
                           n_2818, QN => n1972);
   KEY_EXPAN0_reg_32_9_inst : FD1 port map( D => n5198, CP => CLK_I, Q => 
                           n_2819, QN => n901);
   KEY_EXPAN0_reg_31_9_inst : FD1 port map( D => n5197, CP => CLK_I, Q => 
                           n_2820, QN => n1947);
   KEY_EXPAN0_reg_30_9_inst : FD1 port map( D => n5196, CP => CLK_I, Q => 
                           n_2821, QN => n876);
   KEY_EXPAN0_reg_29_9_inst : FD1 port map( D => n5195, CP => CLK_I, Q => 
                           n_2822, QN => n1946);
   KEY_EXPAN0_reg_28_9_inst : FD1 port map( D => n5194, CP => CLK_I, Q => 
                           n_2823, QN => n875);
   KEY_EXPAN0_reg_27_9_inst : FD1 port map( D => n5193, CP => CLK_I, Q => 
                           n_2824, QN => n1945);
   KEY_EXPAN0_reg_26_9_inst : FD1 port map( D => n5192, CP => CLK_I, Q => 
                           n_2825, QN => n874);
   KEY_EXPAN0_reg_25_9_inst : FD1 port map( D => n5191, CP => CLK_I, Q => 
                           n_2826, QN => n1944);
   KEY_EXPAN0_reg_24_9_inst : FD1 port map( D => n5190, CP => CLK_I, Q => 
                           n_2827, QN => n873);
   KEY_EXPAN0_reg_23_9_inst : FD1 port map( D => n5189, CP => CLK_I, Q => 
                           n_2828, QN => n1951);
   KEY_EXPAN0_reg_22_9_inst : FD1 port map( D => n5188, CP => CLK_I, Q => 
                           n_2829, QN => n880);
   KEY_EXPAN0_reg_21_9_inst : FD1 port map( D => n5187, CP => CLK_I, Q => 
                           n_2830, QN => n1950);
   KEY_EXPAN0_reg_20_9_inst : FD1 port map( D => n5186, CP => CLK_I, Q => 
                           n_2831, QN => n879);
   KEY_EXPAN0_reg_19_9_inst : FD1 port map( D => n5185, CP => CLK_I, Q => 
                           n_2832, QN => n1949);
   KEY_EXPAN0_reg_18_9_inst : FD1 port map( D => n5184, CP => CLK_I, Q => 
                           n_2833, QN => n878);
   KEY_EXPAN0_reg_17_9_inst : FD1 port map( D => n5183, CP => CLK_I, Q => 
                           n_2834, QN => n1948);
   KEY_EXPAN0_reg_16_9_inst : FD1 port map( D => n5182, CP => CLK_I, Q => 
                           n_2835, QN => n877);
   KEY_EXPAN0_reg_15_9_inst : FD1 port map( D => n5181, CP => CLK_I, Q => 
                           n_2836, QN => n1955);
   KEY_EXPAN0_reg_14_9_inst : FD1 port map( D => n5180, CP => CLK_I, Q => 
                           n_2837, QN => n884);
   KEY_EXPAN0_reg_13_9_inst : FD1 port map( D => n5179, CP => CLK_I, Q => 
                           n_2838, QN => n1954);
   KEY_EXPAN0_reg_12_9_inst : FD1 port map( D => n5178, CP => CLK_I, Q => 
                           n_2839, QN => n883);
   KEY_EXPAN0_reg_11_9_inst : FD1 port map( D => n5177, CP => CLK_I, Q => 
                           n_2840, QN => n1953);
   KEY_EXPAN0_reg_10_9_inst : FD1 port map( D => n5176, CP => CLK_I, Q => 
                           n_2841, QN => n882);
   KEY_EXPAN0_reg_9_9_inst : FD1 port map( D => n5175, CP => CLK_I, Q => n_2842
                           , QN => n1952);
   KEY_EXPAN0_reg_8_9_inst : FD1 port map( D => n5174, CP => CLK_I, Q => n_2843
                           , QN => n881);
   KEY_EXPAN0_reg_7_9_inst : FD1 port map( D => n5173, CP => CLK_I, Q => n_2844
                           , QN => n1959);
   KEY_EXPAN0_reg_6_9_inst : FD1 port map( D => n5172, CP => CLK_I, Q => n_2845
                           , QN => n888);
   KEY_EXPAN0_reg_5_9_inst : FD1 port map( D => n5171, CP => CLK_I, Q => n_2846
                           , QN => n1958);
   KEY_EXPAN0_reg_4_9_inst : FD1 port map( D => n5170, CP => CLK_I, Q => n_2847
                           , QN => n887);
   KEY_EXPAN0_reg_3_9_inst : FD1 port map( D => n5169, CP => CLK_I, Q => n_2848
                           , QN => n1957);
   KEY_EXPAN0_reg_2_9_inst : FD1 port map( D => n5168, CP => CLK_I, Q => n_2849
                           , QN => n886);
   KEY_EXPAN0_reg_1_9_inst : FD1 port map( D => n5167, CP => CLK_I, Q => n_2850
                           , QN => n1956);
   KEY_EXPAN0_reg_0_9_inst : FD1 port map( D => n5166, CP => CLK_I, Q => n_2851
                           , QN => n885);
   v_KEY_COL_OUT0_reg_9_inst : FD1 port map( D => n4553, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_9_port, QN => n1045);
   v_TEMP_VECTOR_reg_0_inst : FD1 port map( D => n6695, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_0_port, QN => n_2852);
   KEY_EXPAN0_reg_63_0_inst : FD1 port map( D => n4653, CP => CLK_I, Q => 
                           n_2853, QN => n1995);
   KEY_EXPAN0_reg_62_0_inst : FD1 port map( D => n4652, CP => CLK_I, Q => 
                           n_2854, QN => n924);
   KEY_EXPAN0_reg_61_0_inst : FD1 port map( D => n4651, CP => CLK_I, Q => 
                           n_2855, QN => n1994);
   KEY_EXPAN0_reg_60_0_inst : FD1 port map( D => n4650, CP => CLK_I, Q => 
                           n_2856, QN => n923);
   KEY_EXPAN0_reg_59_0_inst : FD1 port map( D => n4649, CP => CLK_I, Q => 
                           n_2857, QN => n1993);
   KEY_EXPAN0_reg_58_0_inst : FD1 port map( D => n4648, CP => CLK_I, Q => 
                           n_2858, QN => n922);
   KEY_EXPAN0_reg_57_0_inst : FD1 port map( D => n4647, CP => CLK_I, Q => 
                           n_2859, QN => n1992);
   KEY_EXPAN0_reg_56_0_inst : FD1 port map( D => n4646, CP => CLK_I, Q => 
                           n_2860, QN => n921);
   KEY_EXPAN0_reg_55_0_inst : FD1 port map( D => n4645, CP => CLK_I, Q => 
                           n_2861, QN => n1999);
   KEY_EXPAN0_reg_54_0_inst : FD1 port map( D => n4644, CP => CLK_I, Q => 
                           n_2862, QN => n928);
   KEY_EXPAN0_reg_53_0_inst : FD1 port map( D => n4643, CP => CLK_I, Q => 
                           n_2863, QN => n1998);
   KEY_EXPAN0_reg_52_0_inst : FD1 port map( D => n4642, CP => CLK_I, Q => 
                           n_2864, QN => n927);
   KEY_EXPAN0_reg_51_0_inst : FD1 port map( D => n4641, CP => CLK_I, Q => 
                           n_2865, QN => n1997);
   KEY_EXPAN0_reg_50_0_inst : FD1 port map( D => n4640, CP => CLK_I, Q => 
                           n_2866, QN => n926);
   KEY_EXPAN0_reg_49_0_inst : FD1 port map( D => n4639, CP => CLK_I, Q => 
                           n_2867, QN => n1996);
   KEY_EXPAN0_reg_48_0_inst : FD1 port map( D => n4638, CP => CLK_I, Q => 
                           n_2868, QN => n925);
   KEY_EXPAN0_reg_47_0_inst : FD1 port map( D => n4637, CP => CLK_I, Q => 
                           n_2869, QN => n2003);
   KEY_EXPAN0_reg_46_0_inst : FD1 port map( D => n4636, CP => CLK_I, Q => 
                           n_2870, QN => n932);
   KEY_EXPAN0_reg_45_0_inst : FD1 port map( D => n4635, CP => CLK_I, Q => 
                           n_2871, QN => n2002);
   KEY_EXPAN0_reg_44_0_inst : FD1 port map( D => n4634, CP => CLK_I, Q => 
                           n_2872, QN => n931);
   KEY_EXPAN0_reg_43_0_inst : FD1 port map( D => n4633, CP => CLK_I, Q => 
                           n_2873, QN => n2001);
   KEY_EXPAN0_reg_42_0_inst : FD1 port map( D => n4632, CP => CLK_I, Q => 
                           n_2874, QN => n930);
   KEY_EXPAN0_reg_41_0_inst : FD1 port map( D => n4631, CP => CLK_I, Q => 
                           n_2875, QN => n2000);
   KEY_EXPAN0_reg_40_0_inst : FD1 port map( D => n4630, CP => CLK_I, Q => 
                           n_2876, QN => n929);
   KEY_EXPAN0_reg_39_0_inst : FD1 port map( D => n4629, CP => CLK_I, Q => 
                           n_2877, QN => n2007);
   KEY_EXPAN0_reg_38_0_inst : FD1 port map( D => n4628, CP => CLK_I, Q => 
                           n_2878, QN => n936);
   KEY_EXPAN0_reg_37_0_inst : FD1 port map( D => n4627, CP => CLK_I, Q => 
                           n_2879, QN => n2006);
   KEY_EXPAN0_reg_36_0_inst : FD1 port map( D => n4626, CP => CLK_I, Q => 
                           n_2880, QN => n935);
   KEY_EXPAN0_reg_35_0_inst : FD1 port map( D => n4625, CP => CLK_I, Q => 
                           n_2881, QN => n2005);
   KEY_EXPAN0_reg_34_0_inst : FD1 port map( D => n4624, CP => CLK_I, Q => 
                           n_2882, QN => n934);
   KEY_EXPAN0_reg_33_0_inst : FD1 port map( D => n4623, CP => CLK_I, Q => 
                           n_2883, QN => n2004);
   KEY_EXPAN0_reg_32_0_inst : FD1 port map( D => n4622, CP => CLK_I, Q => 
                           n_2884, QN => n933);
   KEY_EXPAN0_reg_31_0_inst : FD1 port map( D => n4621, CP => CLK_I, Q => 
                           n_2885, QN => n1979);
   KEY_EXPAN0_reg_30_0_inst : FD1 port map( D => n4620, CP => CLK_I, Q => 
                           n_2886, QN => n908);
   KEY_EXPAN0_reg_29_0_inst : FD1 port map( D => n4619, CP => CLK_I, Q => 
                           n_2887, QN => n1978);
   KEY_EXPAN0_reg_28_0_inst : FD1 port map( D => n4618, CP => CLK_I, Q => 
                           n_2888, QN => n907);
   KEY_EXPAN0_reg_27_0_inst : FD1 port map( D => n4617, CP => CLK_I, Q => 
                           n_2889, QN => n1977);
   KEY_EXPAN0_reg_26_0_inst : FD1 port map( D => n4616, CP => CLK_I, Q => 
                           n_2890, QN => n906);
   KEY_EXPAN0_reg_25_0_inst : FD1 port map( D => n4615, CP => CLK_I, Q => 
                           n_2891, QN => n1976);
   KEY_EXPAN0_reg_24_0_inst : FD1 port map( D => n4614, CP => CLK_I, Q => 
                           n_2892, QN => n905);
   KEY_EXPAN0_reg_23_0_inst : FD1 port map( D => n4613, CP => CLK_I, Q => 
                           n_2893, QN => n1983);
   KEY_EXPAN0_reg_22_0_inst : FD1 port map( D => n4612, CP => CLK_I, Q => 
                           n_2894, QN => n912);
   KEY_EXPAN0_reg_21_0_inst : FD1 port map( D => n4611, CP => CLK_I, Q => 
                           n_2895, QN => n1982);
   KEY_EXPAN0_reg_20_0_inst : FD1 port map( D => n4610, CP => CLK_I, Q => 
                           n_2896, QN => n911);
   KEY_EXPAN0_reg_19_0_inst : FD1 port map( D => n4609, CP => CLK_I, Q => 
                           n_2897, QN => n1981);
   KEY_EXPAN0_reg_18_0_inst : FD1 port map( D => n4608, CP => CLK_I, Q => 
                           n_2898, QN => n910);
   KEY_EXPAN0_reg_17_0_inst : FD1 port map( D => n4607, CP => CLK_I, Q => 
                           n_2899, QN => n1980);
   KEY_EXPAN0_reg_16_0_inst : FD1 port map( D => n4606, CP => CLK_I, Q => 
                           n_2900, QN => n909);
   KEY_EXPAN0_reg_15_0_inst : FD1 port map( D => n4605, CP => CLK_I, Q => 
                           n_2901, QN => n1987);
   KEY_EXPAN0_reg_14_0_inst : FD1 port map( D => n4604, CP => CLK_I, Q => 
                           n_2902, QN => n916);
   KEY_EXPAN0_reg_13_0_inst : FD1 port map( D => n4603, CP => CLK_I, Q => 
                           n_2903, QN => n1986);
   KEY_EXPAN0_reg_12_0_inst : FD1 port map( D => n4602, CP => CLK_I, Q => 
                           n_2904, QN => n915);
   KEY_EXPAN0_reg_11_0_inst : FD1 port map( D => n4601, CP => CLK_I, Q => 
                           n_2905, QN => n1985);
   KEY_EXPAN0_reg_10_0_inst : FD1 port map( D => n4600, CP => CLK_I, Q => 
                           n_2906, QN => n914);
   KEY_EXPAN0_reg_9_0_inst : FD1 port map( D => n4599, CP => CLK_I, Q => n_2907
                           , QN => n1984);
   KEY_EXPAN0_reg_8_0_inst : FD1 port map( D => n4598, CP => CLK_I, Q => n_2908
                           , QN => n913);
   KEY_EXPAN0_reg_7_0_inst : FD1 port map( D => n4597, CP => CLK_I, Q => n_2909
                           , QN => n1991);
   KEY_EXPAN0_reg_6_0_inst : FD1 port map( D => n4596, CP => CLK_I, Q => n_2910
                           , QN => n920);
   KEY_EXPAN0_reg_5_0_inst : FD1 port map( D => n4595, CP => CLK_I, Q => n_2911
                           , QN => n1990);
   KEY_EXPAN0_reg_4_0_inst : FD1 port map( D => n4594, CP => CLK_I, Q => n_2912
                           , QN => n919);
   KEY_EXPAN0_reg_3_0_inst : FD1 port map( D => n4593, CP => CLK_I, Q => n_2913
                           , QN => n1989);
   KEY_EXPAN0_reg_2_0_inst : FD1 port map( D => n4592, CP => CLK_I, Q => n_2914
                           , QN => n918);
   KEY_EXPAN0_reg_1_0_inst : FD1 port map( D => n4591, CP => CLK_I, Q => n_2915
                           , QN => n1988);
   KEY_EXPAN0_reg_0_0_inst : FD1 port map( D => n4590, CP => CLK_I, Q => n_2916
                           , QN => n917);
   v_KEY_COL_OUT0_reg_0_inst : FD1 port map( D => n4552, CP => CLK_I, Q => 
                           n2110, QN => n4459);
   v_TEMP_VECTOR_reg_24_inst : FD1 port map( D => n6671, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_24_port, QN => n_2917);
   KEY_EXPAN0_reg_63_24_inst : FD1 port map( D => n6189, CP => CLK_I, Q => 
                           n_2918, QN => n2027);
   KEY_EXPAN0_reg_62_24_inst : FD1 port map( D => n6188, CP => CLK_I, Q => 
                           n_2919, QN => n956);
   KEY_EXPAN0_reg_61_24_inst : FD1 port map( D => n6187, CP => CLK_I, Q => 
                           n_2920, QN => n2026);
   KEY_EXPAN0_reg_60_24_inst : FD1 port map( D => n6186, CP => CLK_I, Q => 
                           n_2921, QN => n955);
   KEY_EXPAN0_reg_59_24_inst : FD1 port map( D => n6185, CP => CLK_I, Q => 
                           n_2922, QN => n2025);
   KEY_EXPAN0_reg_58_24_inst : FD1 port map( D => n6184, CP => CLK_I, Q => 
                           n_2923, QN => n954);
   KEY_EXPAN0_reg_57_24_inst : FD1 port map( D => n6183, CP => CLK_I, Q => 
                           n_2924, QN => n2024);
   KEY_EXPAN0_reg_56_24_inst : FD1 port map( D => n6182, CP => CLK_I, Q => 
                           n_2925, QN => n953);
   KEY_EXPAN0_reg_55_24_inst : FD1 port map( D => n6181, CP => CLK_I, Q => 
                           n_2926, QN => n2031);
   KEY_EXPAN0_reg_54_24_inst : FD1 port map( D => n6180, CP => CLK_I, Q => 
                           n_2927, QN => n960);
   KEY_EXPAN0_reg_53_24_inst : FD1 port map( D => n6179, CP => CLK_I, Q => 
                           n_2928, QN => n2030);
   KEY_EXPAN0_reg_52_24_inst : FD1 port map( D => n6178, CP => CLK_I, Q => 
                           n_2929, QN => n959);
   KEY_EXPAN0_reg_51_24_inst : FD1 port map( D => n6177, CP => CLK_I, Q => 
                           n_2930, QN => n2029);
   KEY_EXPAN0_reg_50_24_inst : FD1 port map( D => n6176, CP => CLK_I, Q => 
                           n_2931, QN => n958);
   KEY_EXPAN0_reg_49_24_inst : FD1 port map( D => n6175, CP => CLK_I, Q => 
                           n_2932, QN => n2028);
   KEY_EXPAN0_reg_48_24_inst : FD1 port map( D => n6174, CP => CLK_I, Q => 
                           n_2933, QN => n957);
   KEY_EXPAN0_reg_47_24_inst : FD1 port map( D => n6173, CP => CLK_I, Q => 
                           n_2934, QN => n2035);
   KEY_EXPAN0_reg_46_24_inst : FD1 port map( D => n6172, CP => CLK_I, Q => 
                           n_2935, QN => n964);
   KEY_EXPAN0_reg_45_24_inst : FD1 port map( D => n6171, CP => CLK_I, Q => 
                           n_2936, QN => n2034);
   KEY_EXPAN0_reg_44_24_inst : FD1 port map( D => n6170, CP => CLK_I, Q => 
                           n_2937, QN => n963);
   KEY_EXPAN0_reg_43_24_inst : FD1 port map( D => n6169, CP => CLK_I, Q => 
                           n_2938, QN => n2033);
   KEY_EXPAN0_reg_42_24_inst : FD1 port map( D => n6168, CP => CLK_I, Q => 
                           n_2939, QN => n962);
   KEY_EXPAN0_reg_41_24_inst : FD1 port map( D => n6167, CP => CLK_I, Q => 
                           n_2940, QN => n2032);
   KEY_EXPAN0_reg_40_24_inst : FD1 port map( D => n6166, CP => CLK_I, Q => 
                           n_2941, QN => n961);
   KEY_EXPAN0_reg_39_24_inst : FD1 port map( D => n6165, CP => CLK_I, Q => 
                           n_2942, QN => n2039);
   KEY_EXPAN0_reg_38_24_inst : FD1 port map( D => n6164, CP => CLK_I, Q => 
                           n_2943, QN => n968);
   KEY_EXPAN0_reg_37_24_inst : FD1 port map( D => n6163, CP => CLK_I, Q => 
                           n_2944, QN => n2038);
   KEY_EXPAN0_reg_36_24_inst : FD1 port map( D => n6162, CP => CLK_I, Q => 
                           n_2945, QN => n967);
   KEY_EXPAN0_reg_35_24_inst : FD1 port map( D => n6161, CP => CLK_I, Q => 
                           n_2946, QN => n2037);
   KEY_EXPAN0_reg_34_24_inst : FD1 port map( D => n6160, CP => CLK_I, Q => 
                           n_2947, QN => n966);
   KEY_EXPAN0_reg_33_24_inst : FD1 port map( D => n6159, CP => CLK_I, Q => 
                           n_2948, QN => n2036);
   KEY_EXPAN0_reg_32_24_inst : FD1 port map( D => n6158, CP => CLK_I, Q => 
                           n_2949, QN => n965);
   KEY_EXPAN0_reg_31_24_inst : FD1 port map( D => n6157, CP => CLK_I, Q => 
                           n_2950, QN => n2011);
   KEY_EXPAN0_reg_30_24_inst : FD1 port map( D => n6156, CP => CLK_I, Q => 
                           n_2951, QN => n940);
   KEY_EXPAN0_reg_29_24_inst : FD1 port map( D => n6155, CP => CLK_I, Q => 
                           n_2952, QN => n2010);
   KEY_EXPAN0_reg_28_24_inst : FD1 port map( D => n6154, CP => CLK_I, Q => 
                           n_2953, QN => n939);
   KEY_EXPAN0_reg_27_24_inst : FD1 port map( D => n6153, CP => CLK_I, Q => 
                           n_2954, QN => n2009);
   KEY_EXPAN0_reg_26_24_inst : FD1 port map( D => n6152, CP => CLK_I, Q => 
                           n_2955, QN => n938);
   KEY_EXPAN0_reg_25_24_inst : FD1 port map( D => n6151, CP => CLK_I, Q => 
                           n_2956, QN => n2008);
   KEY_EXPAN0_reg_24_24_inst : FD1 port map( D => n6150, CP => CLK_I, Q => 
                           n_2957, QN => n937);
   KEY_EXPAN0_reg_23_24_inst : FD1 port map( D => n6149, CP => CLK_I, Q => 
                           n_2958, QN => n2015);
   KEY_EXPAN0_reg_22_24_inst : FD1 port map( D => n6148, CP => CLK_I, Q => 
                           n_2959, QN => n944);
   KEY_EXPAN0_reg_21_24_inst : FD1 port map( D => n6147, CP => CLK_I, Q => 
                           n_2960, QN => n2014);
   KEY_EXPAN0_reg_20_24_inst : FD1 port map( D => n6146, CP => CLK_I, Q => 
                           n_2961, QN => n943);
   KEY_EXPAN0_reg_19_24_inst : FD1 port map( D => n6145, CP => CLK_I, Q => 
                           n_2962, QN => n2013);
   KEY_EXPAN0_reg_18_24_inst : FD1 port map( D => n6144, CP => CLK_I, Q => 
                           n_2963, QN => n942);
   KEY_EXPAN0_reg_17_24_inst : FD1 port map( D => n6143, CP => CLK_I, Q => 
                           n_2964, QN => n2012);
   KEY_EXPAN0_reg_16_24_inst : FD1 port map( D => n6142, CP => CLK_I, Q => 
                           n_2965, QN => n941);
   KEY_EXPAN0_reg_15_24_inst : FD1 port map( D => n6141, CP => CLK_I, Q => 
                           n_2966, QN => n2019);
   KEY_EXPAN0_reg_14_24_inst : FD1 port map( D => n6140, CP => CLK_I, Q => 
                           n_2967, QN => n948);
   KEY_EXPAN0_reg_13_24_inst : FD1 port map( D => n6139, CP => CLK_I, Q => 
                           n_2968, QN => n2018);
   KEY_EXPAN0_reg_12_24_inst : FD1 port map( D => n6138, CP => CLK_I, Q => 
                           n_2969, QN => n947);
   KEY_EXPAN0_reg_11_24_inst : FD1 port map( D => n6137, CP => CLK_I, Q => 
                           n_2970, QN => n2017);
   KEY_EXPAN0_reg_10_24_inst : FD1 port map( D => n6136, CP => CLK_I, Q => 
                           n_2971, QN => n946);
   KEY_EXPAN0_reg_9_24_inst : FD1 port map( D => n6135, CP => CLK_I, Q => 
                           n_2972, QN => n2016);
   KEY_EXPAN0_reg_8_24_inst : FD1 port map( D => n6134, CP => CLK_I, Q => 
                           n_2973, QN => n945);
   KEY_EXPAN0_reg_7_24_inst : FD1 port map( D => n6133, CP => CLK_I, Q => 
                           n_2974, QN => n2023);
   KEY_EXPAN0_reg_6_24_inst : FD1 port map( D => n6132, CP => CLK_I, Q => 
                           n_2975, QN => n952);
   KEY_EXPAN0_reg_5_24_inst : FD1 port map( D => n6131, CP => CLK_I, Q => 
                           n_2976, QN => n2022);
   KEY_EXPAN0_reg_4_24_inst : FD1 port map( D => n6130, CP => CLK_I, Q => 
                           n_2977, QN => n951);
   KEY_EXPAN0_reg_3_24_inst : FD1 port map( D => n6129, CP => CLK_I, Q => 
                           n_2978, QN => n2021);
   KEY_EXPAN0_reg_2_24_inst : FD1 port map( D => n6128, CP => CLK_I, Q => 
                           n_2979, QN => n950);
   KEY_EXPAN0_reg_1_24_inst : FD1 port map( D => n6127, CP => CLK_I, Q => 
                           n_2980, QN => n2020);
   KEY_EXPAN0_reg_0_24_inst : FD1 port map( D => n6126, CP => CLK_I, Q => 
                           n_2981, QN => n949);
   v_KEY_COL_OUT0_reg_24_inst : FD1 port map( D => n4551, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_24_port, QN => n1058);
   v_TEMP_VECTOR_reg_16_inst : FD1 port map( D => n6679, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_16_port, QN => n_2982);
   KEY_EXPAN0_reg_63_16_inst : FD1 port map( D => n5677, CP => CLK_I, Q => 
                           n_2983, QN => n2059);
   KEY_EXPAN0_reg_62_16_inst : FD1 port map( D => n5676, CP => CLK_I, Q => 
                           n_2984, QN => n988);
   KEY_EXPAN0_reg_61_16_inst : FD1 port map( D => n5675, CP => CLK_I, Q => 
                           n_2985, QN => n2058);
   KEY_EXPAN0_reg_60_16_inst : FD1 port map( D => n5674, CP => CLK_I, Q => 
                           n_2986, QN => n987);
   KEY_EXPAN0_reg_59_16_inst : FD1 port map( D => n5673, CP => CLK_I, Q => 
                           n_2987, QN => n2057);
   KEY_EXPAN0_reg_58_16_inst : FD1 port map( D => n5672, CP => CLK_I, Q => 
                           n_2988, QN => n986);
   KEY_EXPAN0_reg_57_16_inst : FD1 port map( D => n5671, CP => CLK_I, Q => 
                           n_2989, QN => n2056);
   KEY_EXPAN0_reg_56_16_inst : FD1 port map( D => n5670, CP => CLK_I, Q => 
                           n_2990, QN => n985);
   KEY_EXPAN0_reg_55_16_inst : FD1 port map( D => n5669, CP => CLK_I, Q => 
                           n_2991, QN => n2063);
   KEY_EXPAN0_reg_54_16_inst : FD1 port map( D => n5668, CP => CLK_I, Q => 
                           n_2992, QN => n992);
   KEY_EXPAN0_reg_53_16_inst : FD1 port map( D => n5667, CP => CLK_I, Q => 
                           n_2993, QN => n2062);
   KEY_EXPAN0_reg_52_16_inst : FD1 port map( D => n5666, CP => CLK_I, Q => 
                           n_2994, QN => n991);
   KEY_EXPAN0_reg_51_16_inst : FD1 port map( D => n5665, CP => CLK_I, Q => 
                           n_2995, QN => n2061);
   KEY_EXPAN0_reg_50_16_inst : FD1 port map( D => n5664, CP => CLK_I, Q => 
                           n_2996, QN => n990);
   KEY_EXPAN0_reg_49_16_inst : FD1 port map( D => n5663, CP => CLK_I, Q => 
                           n_2997, QN => n2060);
   KEY_EXPAN0_reg_48_16_inst : FD1 port map( D => n5662, CP => CLK_I, Q => 
                           n_2998, QN => n989);
   KEY_EXPAN0_reg_47_16_inst : FD1 port map( D => n5661, CP => CLK_I, Q => 
                           n_2999, QN => n2067);
   KEY_EXPAN0_reg_46_16_inst : FD1 port map( D => n5660, CP => CLK_I, Q => 
                           n_3000, QN => n996);
   KEY_EXPAN0_reg_45_16_inst : FD1 port map( D => n5659, CP => CLK_I, Q => 
                           n_3001, QN => n2066);
   KEY_EXPAN0_reg_44_16_inst : FD1 port map( D => n5658, CP => CLK_I, Q => 
                           n_3002, QN => n995);
   KEY_EXPAN0_reg_43_16_inst : FD1 port map( D => n5657, CP => CLK_I, Q => 
                           n_3003, QN => n2065);
   KEY_EXPAN0_reg_42_16_inst : FD1 port map( D => n5656, CP => CLK_I, Q => 
                           n_3004, QN => n994);
   KEY_EXPAN0_reg_41_16_inst : FD1 port map( D => n5655, CP => CLK_I, Q => 
                           n_3005, QN => n2064);
   KEY_EXPAN0_reg_40_16_inst : FD1 port map( D => n5654, CP => CLK_I, Q => 
                           n_3006, QN => n993);
   KEY_EXPAN0_reg_39_16_inst : FD1 port map( D => n5653, CP => CLK_I, Q => 
                           n_3007, QN => n2071);
   KEY_EXPAN0_reg_38_16_inst : FD1 port map( D => n5652, CP => CLK_I, Q => 
                           n_3008, QN => n1000);
   KEY_EXPAN0_reg_37_16_inst : FD1 port map( D => n5651, CP => CLK_I, Q => 
                           n_3009, QN => n2070);
   KEY_EXPAN0_reg_36_16_inst : FD1 port map( D => n5650, CP => CLK_I, Q => 
                           n_3010, QN => n999);
   KEY_EXPAN0_reg_35_16_inst : FD1 port map( D => n5649, CP => CLK_I, Q => 
                           n_3011, QN => n2069);
   KEY_EXPAN0_reg_34_16_inst : FD1 port map( D => n5648, CP => CLK_I, Q => 
                           n_3012, QN => n998);
   KEY_EXPAN0_reg_33_16_inst : FD1 port map( D => n5647, CP => CLK_I, Q => 
                           n_3013, QN => n2068);
   KEY_EXPAN0_reg_32_16_inst : FD1 port map( D => n5646, CP => CLK_I, Q => 
                           n_3014, QN => n997);
   KEY_EXPAN0_reg_31_16_inst : FD1 port map( D => n5645, CP => CLK_I, Q => 
                           n_3015, QN => n2043);
   KEY_EXPAN0_reg_30_16_inst : FD1 port map( D => n5644, CP => CLK_I, Q => 
                           n_3016, QN => n972);
   KEY_EXPAN0_reg_29_16_inst : FD1 port map( D => n5643, CP => CLK_I, Q => 
                           n_3017, QN => n2042);
   KEY_EXPAN0_reg_28_16_inst : FD1 port map( D => n5642, CP => CLK_I, Q => 
                           n_3018, QN => n971);
   KEY_EXPAN0_reg_27_16_inst : FD1 port map( D => n5641, CP => CLK_I, Q => 
                           n_3019, QN => n2041);
   KEY_EXPAN0_reg_26_16_inst : FD1 port map( D => n5640, CP => CLK_I, Q => 
                           n_3020, QN => n970);
   KEY_EXPAN0_reg_25_16_inst : FD1 port map( D => n5639, CP => CLK_I, Q => 
                           n_3021, QN => n2040);
   KEY_EXPAN0_reg_24_16_inst : FD1 port map( D => n5638, CP => CLK_I, Q => 
                           n_3022, QN => n969);
   KEY_EXPAN0_reg_23_16_inst : FD1 port map( D => n5637, CP => CLK_I, Q => 
                           n_3023, QN => n2047);
   KEY_EXPAN0_reg_22_16_inst : FD1 port map( D => n5636, CP => CLK_I, Q => 
                           n_3024, QN => n976);
   KEY_EXPAN0_reg_21_16_inst : FD1 port map( D => n5635, CP => CLK_I, Q => 
                           n_3025, QN => n2046);
   KEY_EXPAN0_reg_20_16_inst : FD1 port map( D => n5634, CP => CLK_I, Q => 
                           n_3026, QN => n975);
   KEY_EXPAN0_reg_19_16_inst : FD1 port map( D => n5633, CP => CLK_I, Q => 
                           n_3027, QN => n2045);
   KEY_EXPAN0_reg_18_16_inst : FD1 port map( D => n5632, CP => CLK_I, Q => 
                           n_3028, QN => n974);
   KEY_EXPAN0_reg_17_16_inst : FD1 port map( D => n5631, CP => CLK_I, Q => 
                           n_3029, QN => n2044);
   KEY_EXPAN0_reg_16_16_inst : FD1 port map( D => n5630, CP => CLK_I, Q => 
                           n_3030, QN => n973);
   KEY_EXPAN0_reg_15_16_inst : FD1 port map( D => n5629, CP => CLK_I, Q => 
                           n_3031, QN => n2051);
   KEY_EXPAN0_reg_14_16_inst : FD1 port map( D => n5628, CP => CLK_I, Q => 
                           n_3032, QN => n980);
   KEY_EXPAN0_reg_13_16_inst : FD1 port map( D => n5627, CP => CLK_I, Q => 
                           n_3033, QN => n2050);
   KEY_EXPAN0_reg_12_16_inst : FD1 port map( D => n5626, CP => CLK_I, Q => 
                           n_3034, QN => n979);
   KEY_EXPAN0_reg_11_16_inst : FD1 port map( D => n5625, CP => CLK_I, Q => 
                           n_3035, QN => n2049);
   KEY_EXPAN0_reg_10_16_inst : FD1 port map( D => n5624, CP => CLK_I, Q => 
                           n_3036, QN => n978);
   KEY_EXPAN0_reg_9_16_inst : FD1 port map( D => n5623, CP => CLK_I, Q => 
                           n_3037, QN => n2048);
   KEY_EXPAN0_reg_8_16_inst : FD1 port map( D => n5622, CP => CLK_I, Q => 
                           n_3038, QN => n977);
   KEY_EXPAN0_reg_7_16_inst : FD1 port map( D => n5621, CP => CLK_I, Q => 
                           n_3039, QN => n2055);
   KEY_EXPAN0_reg_6_16_inst : FD1 port map( D => n5620, CP => CLK_I, Q => 
                           n_3040, QN => n984);
   KEY_EXPAN0_reg_5_16_inst : FD1 port map( D => n5619, CP => CLK_I, Q => 
                           n_3041, QN => n2054);
   KEY_EXPAN0_reg_4_16_inst : FD1 port map( D => n5618, CP => CLK_I, Q => 
                           n_3042, QN => n983);
   KEY_EXPAN0_reg_3_16_inst : FD1 port map( D => n5617, CP => CLK_I, Q => 
                           n_3043, QN => n2053);
   KEY_EXPAN0_reg_2_16_inst : FD1 port map( D => n5616, CP => CLK_I, Q => 
                           n_3044, QN => n982);
   KEY_EXPAN0_reg_1_16_inst : FD1 port map( D => n5615, CP => CLK_I, Q => 
                           n_3045, QN => n2052);
   KEY_EXPAN0_reg_0_16_inst : FD1 port map( D => n5614, CP => CLK_I, Q => 
                           n_3046, QN => n981);
   v_KEY_COL_OUT0_reg_16_inst : FD1 port map( D => n4550, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_16_port, QN => n1067);
   v_TEMP_VECTOR_reg_8_inst : FD1 port map( D => n6687, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_8_port, QN => n_3047);
   KEY_EXPAN0_reg_63_8_inst : FD1 port map( D => n5165, CP => CLK_I, Q => 
                           n_3048, QN => n2091);
   KEY_EXPAN0_reg_62_8_inst : FD1 port map( D => n5164, CP => CLK_I, Q => 
                           n_3049, QN => n1020);
   KEY_EXPAN0_reg_61_8_inst : FD1 port map( D => n5163, CP => CLK_I, Q => 
                           n_3050, QN => n2090);
   KEY_EXPAN0_reg_60_8_inst : FD1 port map( D => n5162, CP => CLK_I, Q => 
                           n_3051, QN => n1019);
   KEY_EXPAN0_reg_59_8_inst : FD1 port map( D => n5161, CP => CLK_I, Q => 
                           n_3052, QN => n2089);
   KEY_EXPAN0_reg_58_8_inst : FD1 port map( D => n5160, CP => CLK_I, Q => 
                           n_3053, QN => n1018);
   KEY_EXPAN0_reg_57_8_inst : FD1 port map( D => n5159, CP => CLK_I, Q => 
                           n_3054, QN => n2088);
   KEY_EXPAN0_reg_56_8_inst : FD1 port map( D => n5158, CP => CLK_I, Q => 
                           n_3055, QN => n1017);
   KEY_EXPAN0_reg_55_8_inst : FD1 port map( D => n5157, CP => CLK_I, Q => 
                           n_3056, QN => n2095);
   KEY_EXPAN0_reg_54_8_inst : FD1 port map( D => n5156, CP => CLK_I, Q => 
                           n_3057, QN => n1024);
   KEY_EXPAN0_reg_53_8_inst : FD1 port map( D => n5155, CP => CLK_I, Q => 
                           n_3058, QN => n2094);
   KEY_EXPAN0_reg_52_8_inst : FD1 port map( D => n5154, CP => CLK_I, Q => 
                           n_3059, QN => n1023);
   KEY_EXPAN0_reg_51_8_inst : FD1 port map( D => n5153, CP => CLK_I, Q => 
                           n_3060, QN => n2093);
   KEY_EXPAN0_reg_50_8_inst : FD1 port map( D => n5152, CP => CLK_I, Q => 
                           n_3061, QN => n1022);
   KEY_EXPAN0_reg_49_8_inst : FD1 port map( D => n5151, CP => CLK_I, Q => 
                           n_3062, QN => n2092);
   KEY_EXPAN0_reg_48_8_inst : FD1 port map( D => n5150, CP => CLK_I, Q => 
                           n_3063, QN => n1021);
   KEY_EXPAN0_reg_47_8_inst : FD1 port map( D => n5149, CP => CLK_I, Q => 
                           n_3064, QN => n2099);
   KEY_EXPAN0_reg_46_8_inst : FD1 port map( D => n5148, CP => CLK_I, Q => 
                           n_3065, QN => n1028);
   KEY_EXPAN0_reg_45_8_inst : FD1 port map( D => n5147, CP => CLK_I, Q => 
                           n_3066, QN => n2098);
   KEY_EXPAN0_reg_44_8_inst : FD1 port map( D => n5146, CP => CLK_I, Q => 
                           n_3067, QN => n1027);
   KEY_EXPAN0_reg_43_8_inst : FD1 port map( D => n5145, CP => CLK_I, Q => 
                           n_3068, QN => n2097);
   KEY_EXPAN0_reg_42_8_inst : FD1 port map( D => n5144, CP => CLK_I, Q => 
                           n_3069, QN => n1026);
   KEY_EXPAN0_reg_41_8_inst : FD1 port map( D => n5143, CP => CLK_I, Q => 
                           n_3070, QN => n2096);
   KEY_EXPAN0_reg_40_8_inst : FD1 port map( D => n5142, CP => CLK_I, Q => 
                           n_3071, QN => n1025);
   KEY_EXPAN0_reg_39_8_inst : FD1 port map( D => n5141, CP => CLK_I, Q => 
                           n_3072, QN => n2103);
   KEY_EXPAN0_reg_38_8_inst : FD1 port map( D => n5140, CP => CLK_I, Q => 
                           n_3073, QN => n1032);
   KEY_EXPAN0_reg_37_8_inst : FD1 port map( D => n5139, CP => CLK_I, Q => 
                           n_3074, QN => n2102);
   KEY_EXPAN0_reg_36_8_inst : FD1 port map( D => n5138, CP => CLK_I, Q => 
                           n_3075, QN => n1031);
   KEY_EXPAN0_reg_35_8_inst : FD1 port map( D => n5137, CP => CLK_I, Q => 
                           n_3076, QN => n2101);
   KEY_EXPAN0_reg_34_8_inst : FD1 port map( D => n5136, CP => CLK_I, Q => 
                           n_3077, QN => n1030);
   KEY_EXPAN0_reg_33_8_inst : FD1 port map( D => n5135, CP => CLK_I, Q => 
                           n_3078, QN => n2100);
   KEY_EXPAN0_reg_32_8_inst : FD1 port map( D => n5134, CP => CLK_I, Q => 
                           n_3079, QN => n1029);
   KEY_EXPAN0_reg_31_8_inst : FD1 port map( D => n5133, CP => CLK_I, Q => 
                           n_3080, QN => n2075);
   KEY_EXPAN0_reg_30_8_inst : FD1 port map( D => n5132, CP => CLK_I, Q => 
                           n_3081, QN => n1004);
   KEY_EXPAN0_reg_29_8_inst : FD1 port map( D => n5131, CP => CLK_I, Q => 
                           n_3082, QN => n2074);
   KEY_EXPAN0_reg_28_8_inst : FD1 port map( D => n5130, CP => CLK_I, Q => 
                           n_3083, QN => n1003);
   KEY_EXPAN0_reg_27_8_inst : FD1 port map( D => n5129, CP => CLK_I, Q => 
                           n_3084, QN => n2073);
   KEY_EXPAN0_reg_26_8_inst : FD1 port map( D => n5128, CP => CLK_I, Q => 
                           n_3085, QN => n1002);
   KEY_EXPAN0_reg_25_8_inst : FD1 port map( D => n5127, CP => CLK_I, Q => 
                           n_3086, QN => n2072);
   KEY_EXPAN0_reg_24_8_inst : FD1 port map( D => n5126, CP => CLK_I, Q => 
                           n_3087, QN => n1001);
   KEY_EXPAN0_reg_23_8_inst : FD1 port map( D => n5125, CP => CLK_I, Q => 
                           n_3088, QN => n2079);
   KEY_EXPAN0_reg_22_8_inst : FD1 port map( D => n5124, CP => CLK_I, Q => 
                           n_3089, QN => n1008);
   KEY_EXPAN0_reg_21_8_inst : FD1 port map( D => n5123, CP => CLK_I, Q => 
                           n_3090, QN => n2078);
   KEY_EXPAN0_reg_20_8_inst : FD1 port map( D => n5122, CP => CLK_I, Q => 
                           n_3091, QN => n1007);
   KEY_EXPAN0_reg_19_8_inst : FD1 port map( D => n5121, CP => CLK_I, Q => 
                           n_3092, QN => n2077);
   KEY_EXPAN0_reg_18_8_inst : FD1 port map( D => n5120, CP => CLK_I, Q => 
                           n_3093, QN => n1006);
   KEY_EXPAN0_reg_17_8_inst : FD1 port map( D => n5119, CP => CLK_I, Q => 
                           n_3094, QN => n2076);
   KEY_EXPAN0_reg_16_8_inst : FD1 port map( D => n5118, CP => CLK_I, Q => 
                           n_3095, QN => n1005);
   KEY_EXPAN0_reg_15_8_inst : FD1 port map( D => n5117, CP => CLK_I, Q => 
                           n_3096, QN => n2083);
   KEY_EXPAN0_reg_14_8_inst : FD1 port map( D => n5116, CP => CLK_I, Q => 
                           n_3097, QN => n1012);
   KEY_EXPAN0_reg_13_8_inst : FD1 port map( D => n5115, CP => CLK_I, Q => 
                           n_3098, QN => n2082);
   KEY_EXPAN0_reg_12_8_inst : FD1 port map( D => n5114, CP => CLK_I, Q => 
                           n_3099, QN => n1011);
   KEY_EXPAN0_reg_11_8_inst : FD1 port map( D => n5113, CP => CLK_I, Q => 
                           n_3100, QN => n2081);
   KEY_EXPAN0_reg_10_8_inst : FD1 port map( D => n5112, CP => CLK_I, Q => 
                           n_3101, QN => n1010);
   KEY_EXPAN0_reg_9_8_inst : FD1 port map( D => n5111, CP => CLK_I, Q => n_3102
                           , QN => n2080);
   KEY_EXPAN0_reg_8_8_inst : FD1 port map( D => n5110, CP => CLK_I, Q => n_3103
                           , QN => n1009);
   KEY_EXPAN0_reg_7_8_inst : FD1 port map( D => n5109, CP => CLK_I, Q => n_3104
                           , QN => n2087);
   KEY_EXPAN0_reg_6_8_inst : FD1 port map( D => n5108, CP => CLK_I, Q => n_3105
                           , QN => n1016);
   KEY_EXPAN0_reg_5_8_inst : FD1 port map( D => n5107, CP => CLK_I, Q => n_3106
                           , QN => n2086);
   KEY_EXPAN0_reg_4_8_inst : FD1 port map( D => n5106, CP => CLK_I, Q => n_3107
                           , QN => n1015);
   KEY_EXPAN0_reg_3_8_inst : FD1 port map( D => n5105, CP => CLK_I, Q => n_3108
                           , QN => n2085);
   KEY_EXPAN0_reg_2_8_inst : FD1 port map( D => n5104, CP => CLK_I, Q => n_3109
                           , QN => n1014);
   KEY_EXPAN0_reg_1_8_inst : FD1 port map( D => n5103, CP => CLK_I, Q => n_3110
                           , QN => n2084);
   KEY_EXPAN0_reg_0_8_inst : FD1 port map( D => n5102, CP => CLK_I, Q => n_3111
                           , QN => n1013);
   v_KEY_COL_OUT0_reg_8_inst : FD1 port map( D => n4549, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_8_port, QN => n1046);
   U3 : MUX21H port map( A => v_KEY32_IN_24_port, B => KEY_I(0), S => n2121, Z 
                           => n4472);
   U4 : MUX21H port map( A => v_KEY32_IN_25_port, B => KEY_I(1), S => n2121, Z 
                           => n4473);
   U5 : MUX21H port map( A => v_KEY32_IN_26_port, B => KEY_I(2), S => n2121, Z 
                           => n4474);
   U6 : MUX21H port map( A => v_KEY32_IN_27_port, B => KEY_I(3), S => n2121, Z 
                           => n4475);
   U7 : MUX21H port map( A => v_KEY32_IN_28_port, B => KEY_I(4), S => n2121, Z 
                           => n4476);
   U8 : MUX21H port map( A => v_KEY32_IN_29_port, B => KEY_I(5), S => n2121, Z 
                           => n4477);
   U9 : MUX21H port map( A => v_KEY32_IN_30_port, B => KEY_I(6), S => n2121, Z 
                           => n4478);
   U10 : MUX21H port map( A => v_KEY32_IN_31_port, B => KEY_I(7), S => n2121, Z
                           => n4479);
   U11 : MUX21H port map( A => v_KEY32_IN_0_port, B => KEY_I(0), S => n2122, Z 
                           => n4480);
   U12 : MUX21H port map( A => v_KEY32_IN_1_port, B => KEY_I(1), S => n2122, Z 
                           => n4481);
   U13 : MUX21H port map( A => v_KEY32_IN_2_port, B => KEY_I(2), S => n2122, Z 
                           => n4482);
   U14 : MUX21H port map( A => v_KEY32_IN_3_port, B => KEY_I(3), S => n2122, Z 
                           => n4483);
   U15 : MUX21H port map( A => v_KEY32_IN_4_port, B => KEY_I(4), S => n2122, Z 
                           => n4484);
   U16 : MUX21H port map( A => v_KEY32_IN_5_port, B => KEY_I(5), S => n2122, Z 
                           => n4485);
   U17 : MUX21H port map( A => v_KEY32_IN_6_port, B => KEY_I(6), S => n2122, Z 
                           => n4486);
   U18 : MUX21H port map( A => v_KEY32_IN_7_port, B => KEY_I(7), S => n2122, Z 
                           => n4487);
   U19 : AN3 port map( A => n6, B => n1039, C => n2123, Z => n2122);
   U20 : MUX21H port map( A => v_KEY32_IN_16_port, B => KEY_I(0), S => n2124, Z
                           => n4488);
   U21 : MUX21H port map( A => v_KEY32_IN_17_port, B => KEY_I(1), S => n2124, Z
                           => n4489);
   U22 : MUX21H port map( A => v_KEY32_IN_18_port, B => KEY_I(2), S => n2124, Z
                           => n4490);
   U23 : MUX21H port map( A => v_KEY32_IN_19_port, B => KEY_I(3), S => n2124, Z
                           => n4491);
   U24 : MUX21H port map( A => v_KEY32_IN_20_port, B => KEY_I(4), S => n2124, Z
                           => n4492);
   U25 : MUX21H port map( A => v_KEY32_IN_21_port, B => KEY_I(5), S => n2124, Z
                           => n4493);
   U26 : MUX21H port map( A => v_KEY32_IN_22_port, B => KEY_I(6), S => n2124, Z
                           => n4494);
   U27 : MUX21H port map( A => v_KEY32_IN_23_port, B => KEY_I(7), S => n2124, Z
                           => n4495);
   U28 : AN3 port map( A => n1039, B => n2123, C => n4463, Z => n2124);
   U29 : MUX21H port map( A => KEY_I(0), B => v_KEY32_IN_8_port, S => n2125, Z 
                           => n4496);
   U30 : MUX21H port map( A => KEY_I(1), B => v_KEY32_IN_9_port, S => n2125, Z 
                           => n4497);
   U31 : MUX21H port map( A => KEY_I(2), B => v_KEY32_IN_10_port, S => n2125, Z
                           => n4498);
   U32 : MUX21H port map( A => KEY_I(3), B => v_KEY32_IN_11_port, S => n2125, Z
                           => n4499);
   U33 : MUX21H port map( A => KEY_I(4), B => v_KEY32_IN_12_port, S => n2125, Z
                           => n4500);
   U34 : MUX21H port map( A => KEY_I(5), B => v_KEY32_IN_13_port, S => n2125, Z
                           => n4501);
   U35 : MUX21H port map( A => KEY_I(6), B => v_KEY32_IN_14_port, S => n2125, Z
                           => n4502);
   U36 : MUX21H port map( A => KEY_I(7), B => v_KEY32_IN_15_port, S => n2125, Z
                           => n4503);
   U37 : MUX21L port map( A => n2126, B => n2127, S => 
                           v_CALCULATION_CNTR_5_port, Z => n4504);
   U38 : ND2 port map( A => n2128, B => n2129, Z => n2126);
   U39 : MUX21H port map( A => n2130, B => n2131, S => n1079, Z => n4505);
   U40 : MUX21L port map( A => n2132, B => n2133, S => 
                           v_CALCULATION_CNTR_7_port, Z => n4506);
   U41 : AO6 port map( A => n2128, B => n1079, C => n2130, Z => n2133);
   U42 : AO7 port map( A => v_CALCULATION_CNTR_5_port, B => n2134, C => n2127, 
                           Z => n2130);
   U43 : IV port map( A => n2135, Z => n2127);
   U44 : AO7 port map( A => n2129, B => n2134, C => n2136, Z => n2135);
   U45 : ND2 port map( A => n2131, B => v_CALCULATION_CNTR_6_port, Z => n2132);
   U46 : AN3 port map( A => n2128, B => n2129, C => v_CALCULATION_CNTR_5_port, 
                           Z => n2131);
   U47 : NR3 port map( A => n2137, B => n8, C => n1078, Z => n2129);
   U48 : MUX21L port map( A => n2138, B => CE_I, S => n4464, Z => n6749);
   U49 : AO7 port map( A => n2139, B => n6, C => n2125, Z => n6748);
   U50 : ND3 port map( A => n6, B => n2123, C => n4464, Z => n2125);
   U51 : AO6 port map( A => VALID_KEY_I, B => n1039, C => n2140, Z => n2139);
   U52 : MUX21L port map( A => n2141, B => n2142, S => n4462, Z => n6715);
   U53 : AO6 port map( A => n2143, B => n2144, C => n2145, Z => n2142);
   U54 : IV port map( A => n2146, Z => n2144);
   U55 : ND2 port map( A => n2146, B => n2147, Z => n2141);
   U56 : MUX21H port map( A => n2145, B => n2147, S => n3, Z => n6714);
   U57 : MUX21L port map( A => n2148, B => n2149, S => n4460, Z => n6713);
   U58 : ND2 port map( A => n2147, B => n4461, Z => n2148);
   U59 : AO7 port map( A => n2149, B => n5, C => n2150, Z => n6712);
   U60 : AO2 port map( A => n2151, B => n2143, C => n2152, D => n2147, Z => 
                           n2150);
   U61 : NR2 port map( A => n2145, B => n2153, Z => n2147);
   U62 : AO6 port map( A => n3, B => n2143, C => n2145, Z => n2149);
   U63 : AO7 port map( A => n2154, B => n2155, C => n2156, Z => n2145);
   U64 : MUX21L port map( A => n2157, B => n1043, S => n2158, Z => n6711);
   U65 : NR2 port map( A => n2159, B => n2160, Z => n2158);
   U66 : AO6 port map( A => n2146, B => n1042, C => n2140, Z => n2159);
   U67 : MUX21L port map( A => n2161, B => n2489, S => n2162, Z => n6710);
   U68 : ND2 port map( A => n2163, B => n2164, Z => n2161);
   U69 : MUX21L port map( A => n2157, B => n4455, S => n2162, Z => n6709);
   U70 : NR2 port map( A => n2160, B => n2165, Z => n2162);
   U71 : AN3 port map( A => CE_I, B => n1042, C => n2146, Z => n2165);
   U72 : AO7 port map( A => n2140, B => n2163, C => n2164, Z => n2160);
   U73 : IV port map( A => n2166, Z => n2163);
   U74 : ND2 port map( A => n2166, B => n2164, Z => n2157);
   U75 : NR2 port map( A => n1040, B => VALID_KEY_I, Z => n2166);
   U76 : MUX21L port map( A => n2167, B => n2168, S => n6649, Z => n6708);
   U77 : MUX21L port map( A => n2169, B => n2170, S => n6648, Z => n6707);
   U78 : ND2 port map( A => n2171, B => n1, Z => n2170);
   U79 : IV port map( A => n2172, Z => n2169);
   U80 : MUX21L port map( A => n2173, B => n2174, S => n6647, Z => n6706);
   U81 : ND3 port map( A => n1033, B => n1, C => n2171, Z => n2174);
   U82 : AO6 port map( A => n6648, B => n2171, C => n2172, Z => n2173);
   U83 : AO7 port map( A => n2168, B => n1, C => n2167, Z => n2172);
   U84 : MUX21L port map( A => n2175, B => n2176, S => n6646, Z => n6705);
   U85 : ND2 port map( A => n2177, B => n2171, Z => n2176);
   U86 : MUX21H port map( A => n2178, B => n2179, S => n1037, Z => n6704);
   U87 : MUX21L port map( A => n2180, B => n2181, S => n6644, Z => n6703);
   U88 : ND2 port map( A => n2178, B => n1037, Z => n2181);
   U89 : AN3 port map( A => n2171, B => n1044, C => n2177, Z => n2178);
   U90 : AO6 port map( A => n6645, B => n2171, C => n2179, Z => n2180);
   U91 : AO7 port map( A => n2168, B => n1044, C => n2175, Z => n2179);
   U92 : IV port map( A => n2182, Z => n2175);
   U93 : AO7 port map( A => n2177, B => n2168, C => n2167, Z => n2182);
   U94 : NR3 port map( A => n6649, B => n6648, C => n6647, Z => n2177);
   U95 : IV port map( A => n2168, Z => n2171);
   U96 : ND2 port map( A => n2183, B => n2167, Z => n2168);
   U97 : AO7 port map( A => n2184, B => n2140, C => n2185, Z => n2167);
   U98 : AO6 port map( A => n2186, B => n1036, C => n2187, Z => n2184);
   U99 : AO7 port map( A => n2188, B => n2189, C => n2190, Z => n2186);
   U100 : AO4 port map( A => n2136, B => n1076, C => RESET_I, D => n2191, Z => 
                           n6702);
   U101 : AO6 port map( A => CE_I, B => n2192, C => n2121, Z => n2191);
   U102 : AN3 port map( A => n2123, B => n4464, C => n4463, Z => n2121);
   U103 : MUX21L port map( A => n2193, B => n2194, S => n6638, Z => n6701);
   U104 : ND2 port map( A => n2195, B => n2, Z => n2194);
   U105 : AO6 port map( A => n6639, B => n2196, C => n2197, Z => n2193);
   U106 : MUX21L port map( A => n2198, B => n2199, S => n6643, Z => n6700);
   U107 : EON1 port map( A => n2199, B => n2200, C => n1038, D => n2201, Z => 
                           n6699);
   U108 : AO4 port map( A => n2199, B => n2202, C => n6641, D => n2203, Z => 
                           n6698);
   U109 : AO6 port map( A => n6642, B => n2196, C => n2201, Z => n2203);
   U110 : AO7 port map( A => n2199, B => n4, C => n2198, Z => n2201);
   U111 : MUX21L port map( A => n2204, B => n2205, S => n6640, Z => n6697);
   U112 : ND2 port map( A => n2206, B => n2196, Z => n2205);
   U113 : MUX21H port map( A => n2195, B => n2197, S => n2, Z => n6696);
   U114 : AO7 port map( A => n2199, B => n1035, C => n2204, Z => n2197);
   U115 : IV port map( A => n2207, Z => n2204);
   U116 : AO7 port map( A => n2206, B => n2199, C => n2198, Z => n2207);
   U117 : AN3 port map( A => n2196, B => n1035, C => n2206, Z => n2195);
   U118 : IV port map( A => n2199, Z => n2196);
   U119 : ND2 port map( A => n2183, B => n2198, Z => n2199);
   U120 : AO7 port map( A => n2140, B => n1076, C => n2185, Z => n2198);
   U121 : AO6 port map( A => n1040, B => n2123, C => RESET_I, Z => n2185);
   U122 : IV port map( A => n2138, Z => n2123);
   U123 : AO6 port map( A => n1040, B => VALID_KEY_I, C => RESET_I, Z => n2183)
                           ;
   U124 : AO3 port map( A => n2109, B => n2208, C => n2209, D => n2210, Z => 
                           n6695);
   U125 : AO2 port map( A => n2211, B => n2212, C => v_SUB_WORD_0_port, D => 
                           n2213, Z => n2210);
   U126 : EN port map( A => n2214, B => v_TEMP_VECTOR_8_port, Z => n2212);
   U127 : OR3 port map( A => n4458, B => n4460, C => n4461, Z => n2214);
   U128 : MUX21L port map( A => n2215, B => n2216, S => v_TEMP_VECTOR_0_port, Z
                           => n2209);
   U129 : AO7 port map( A => n2217, B => n2110, C => n2218, Z => n2216);
   U130 : NR2 port map( A => n4459, B => n2217, Z => n2215);
   U131 : AO3 port map( A => n2111, B => n2208, C => n2219, D => n2220, Z => 
                           n6694);
   U132 : AO2 port map( A => n2221, B => n2211, C => n2213, D => n2108, Z => 
                           n2220);
   U133 : EN port map( A => n2222, B => v_TEMP_VECTOR_9_port, Z => n2221);
   U134 : AO6 port map( A => n2223, B => n4461, C => n4462, Z => n2222);
   U135 : NR2 port map( A => n4458, B => n4460, Z => n2223);
   U136 : MUX21L port map( A => n2224, B => n2225, S => v_TEMP_VECTOR_1_port, Z
                           => n2219);
   U137 : AO7 port map( A => v_KEY_COL_OUT0_1_port, B => n2217, C => n2218, Z 
                           => n2225);
   U138 : NR2 port map( A => n2217, B => n1063, Z => n2224);
   U139 : AO3 port map( A => n2112, B => n2208, C => n2226, D => n2227, Z => 
                           n6693);
   U140 : AO2 port map( A => n2211, B => n2228, C => n2213, D => n2113, Z => 
                           n2227);
   U141 : EO port map( A => v_TEMP_VECTOR_10_port, B => n2229, Z => n2228);
   U142 : MUX21L port map( A => n2230, B => n1042, S => n4461, Z => n2229);
   U143 : ND2 port map( A => n4460, B => n5, Z => n2230);
   U144 : MUX21L port map( A => n2231, B => n2232, S => v_TEMP_VECTOR_2_port, Z
                           => n2226);
   U145 : AO7 port map( A => v_KEY_COL_OUT0_2_port, B => n2217, C => n2218, Z 
                           => n2232);
   U146 : NR2 port map( A => n2217, B => n1052, Z => n2231);
   U147 : AO3 port map( A => n2114, B => n2208, C => n2233, D => n2234, Z => 
                           n6692);
   U148 : AO2 port map( A => n2235, B => n2211, C => n2213, D => n2107, Z => 
                           n2234);
   U149 : EN port map( A => n2236, B => v_TEMP_VECTOR_11_port, Z => n2235);
   U150 : AO6 port map( A => n4462, B => n3, C => n2152, Z => n2236);
   U151 : NR3 port map( A => n3, B => n4458, C => n2104, Z => n2152);
   U152 : MUX21L port map( A => n2237, B => n2238, S => v_TEMP_VECTOR_3_port, Z
                           => n2233);
   U153 : AO7 port map( A => v_KEY_COL_OUT0_3_port, B => n2217, C => n2218, Z 
                           => n2238);
   U154 : NR2 port map( A => n2217, B => n1049, Z => n2237);
   U155 : AO3 port map( A => n2115, B => n2208, C => n2239, D => n2240, Z => 
                           n6691);
   U156 : AO2 port map( A => n2241, B => n2211, C => n2213, D => n2106, Z => 
                           n2240);
   U157 : EN port map( A => v_TEMP_VECTOR_12_port, B => n2242, Z => n2241);
   U158 : AO6 port map( A => n3, B => n2151, C => n4462, Z => n2242);
   U159 : MUX21L port map( A => n2243, B => n2244, S => v_TEMP_VECTOR_4_port, Z
                           => n2239);
   U160 : AO7 port map( A => v_KEY_COL_OUT0_4_port, B => n2217, C => n2218, Z 
                           => n2244);
   U161 : NR2 port map( A => n2217, B => n1048, Z => n2243);
   U162 : AO3 port map( A => n2116, B => n2208, C => n2245, D => n2246, Z => 
                           n6690);
   U163 : AO2 port map( A => n2211, B => n2247, C => n2213, D => n2105, Z => 
                           n2246);
   U164 : EN port map( A => n2248, B => v_TEMP_VECTOR_13_port, Z => n2247);
   U165 : AO7 port map( A => n2151, B => n4462, C => n4461, Z => n2248);
   U166 : NR2 port map( A => n5, B => n4460, Z => n2151);
   U167 : MUX21L port map( A => n2249, B => n2250, S => v_TEMP_VECTOR_5_port, Z
                           => n2245);
   U168 : AO7 port map( A => v_KEY_COL_OUT0_5_port, B => n2217, C => n2218, Z 
                           => n2250);
   U169 : NR2 port map( A => n2217, B => n1047, Z => n2249);
   U170 : AO3 port map( A => n2117, B => n2208, C => n2251, D => n2252, Z => 
                           n6689);
   U171 : AO2 port map( A => n2211, B => n2253, C => v_SUB_WORD_6_port, D => 
                           n2213, Z => n2252);
   U172 : EN port map( A => n2254, B => v_TEMP_VECTOR_14_port, Z => n2253);
   U173 : OR3 port map( A => n4461, B => n2104, C => n5, Z => n2254);
   U174 : MUX21L port map( A => n2255, B => n2256, S => v_TEMP_VECTOR_6_port, Z
                           => n2251);
   U175 : AO7 port map( A => n2217, B => n2118, C => n2218, Z => n2256);
   U176 : NR2 port map( A => n4457, B => n2217, Z => n2255);
   U177 : AO3 port map( A => n2119, B => n2208, C => n2257, D => n2258, Z => 
                           n6688);
   U178 : AO2 port map( A => n2211, B => n2259, C => v_SUB_WORD_7_port, D => 
                           n2213, Z => n2258);
   U179 : NR2 port map( A => n2260, B => n2261, Z => n2213);
   U180 : EO port map( A => n2146, B => v_TEMP_VECTOR_15_port, Z => n2259);
   U181 : AN3 port map( A => n4460, B => n4461, C => n4458, Z => n2146);
   U182 : NR2 port map( A => n2260, B => n2262, Z => n2211);
   U183 : MUX21L port map( A => n2263, B => n2264, S => v_TEMP_VECTOR_7_port, Z
                           => n2257);
   U184 : AO7 port map( A => n2217, B => n2120, C => n2218, Z => n2264);
   U185 : NR2 port map( A => n4454, B => n2217, Z => n2263);
   U186 : OR2 port map( A => n2260, B => n2265, Z => n2217);
   U187 : ND2 port map( A => n2143, B => n2218, Z => n2260);
   U188 : ND2 port map( A => n2266, B => n2218, Z => n2208);
   U189 : ND2 port map( A => n2267, B => n2268, Z => n2218);
   U190 : AO7 port map( A => n2265, B => n2192, C => CE_I, Z => n2268);
   U191 : ND2 port map( A => n2261, B => n2262, Z => n2265);
   U192 : AO3 port map( A => n1074, B => n2269, C => n2270, D => n2271, Z => 
                           n6687);
   U193 : AO2 port map( A => n2272, B => v_KEY32_IN_8_port, C => 
                           v_TEMP_VECTOR_16_port, D => n2273, Z => n2271);
   U194 : MUX21L port map( A => n2274, B => n2275, S => v_TEMP_VECTOR_8_port, Z
                           => n2270);
   U195 : AO7 port map( A => v_KEY_COL_OUT0_8_port, B => n2276, C => n2277, Z 
                           => n2275);
   U196 : NR2 port map( A => n2276, B => n1046, Z => n2274);
   U197 : AO3 port map( A => n4456, B => n2269, C => n2278, D => n2279, Z => 
                           n6686);
   U198 : AO2 port map( A => n2272, B => v_KEY32_IN_9_port, C => 
                           v_TEMP_VECTOR_17_port, D => n2273, Z => n2279);
   U199 : MUX21L port map( A => n2280, B => n2281, S => v_TEMP_VECTOR_9_port, Z
                           => n2278);
   U200 : AO7 port map( A => v_KEY_COL_OUT0_9_port, B => n2276, C => n2277, Z 
                           => n2281);
   U201 : NR2 port map( A => n2276, B => n1045, Z => n2280);
   U202 : AO3 port map( A => n4465, B => n2269, C => n2282, D => n2283, Z => 
                           n6685);
   U203 : AO2 port map( A => n2272, B => v_KEY32_IN_10_port, C => 
                           v_TEMP_VECTOR_18_port, D => n2273, Z => n2283);
   U204 : MUX21L port map( A => n2284, B => n2285, S => v_TEMP_VECTOR_10_port, 
                           Z => n2282);
   U205 : AO7 port map( A => v_KEY_COL_OUT0_10_port, B => n2276, C => n2277, Z 
                           => n2285);
   U206 : NR2 port map( A => n2276, B => n1073, Z => n2284);
   U207 : AO3 port map( A => n4466, B => n2269, C => n2286, D => n2287, Z => 
                           n6684);
   U208 : AO2 port map( A => n2272, B => v_KEY32_IN_11_port, C => 
                           v_TEMP_VECTOR_19_port, D => n2273, Z => n2287);
   U209 : MUX21L port map( A => n2288, B => n2289, S => v_TEMP_VECTOR_11_port, 
                           Z => n2286);
   U210 : AO7 port map( A => v_KEY_COL_OUT0_11_port, B => n2276, C => n2277, Z 
                           => n2289);
   U211 : NR2 port map( A => n2276, B => n1072, Z => n2288);
   U212 : AO3 port map( A => n4467, B => n2269, C => n2290, D => n2291, Z => 
                           n6683);
   U213 : AO2 port map( A => n2272, B => v_KEY32_IN_12_port, C => 
                           v_TEMP_VECTOR_20_port, D => n2273, Z => n2291);
   U214 : MUX21L port map( A => n2292, B => n2293, S => v_TEMP_VECTOR_12_port, 
                           Z => n2290);
   U215 : AO7 port map( A => v_KEY_COL_OUT0_12_port, B => n2276, C => n2277, Z 
                           => n2293);
   U216 : NR2 port map( A => n2276, B => n1071, Z => n2292);
   U217 : AO3 port map( A => n4468, B => n2269, C => n2294, D => n2295, Z => 
                           n6682);
   U218 : AO2 port map( A => n2272, B => v_KEY32_IN_13_port, C => 
                           v_TEMP_VECTOR_21_port, D => n2273, Z => n2295);
   U219 : MUX21L port map( A => n2296, B => n2297, S => v_TEMP_VECTOR_13_port, 
                           Z => n2294);
   U220 : AO7 port map( A => v_KEY_COL_OUT0_13_port, B => n2276, C => n2277, Z 
                           => n2297);
   U221 : NR2 port map( A => n2276, B => n1070, Z => n2296);
   U222 : AO3 port map( A => n1041, B => n2269, C => n2298, D => n2299, Z => 
                           n6681);
   U223 : AO2 port map( A => n2272, B => v_KEY32_IN_14_port, C => 
                           v_TEMP_VECTOR_22_port, D => n2273, Z => n2299);
   U224 : MUX21L port map( A => n2300, B => n2301, S => v_TEMP_VECTOR_14_port, 
                           Z => n2298);
   U225 : AO7 port map( A => v_KEY_COL_OUT0_14_port, B => n2276, C => n2277, Z 
                           => n2301);
   U226 : NR2 port map( A => n2276, B => n1069, Z => n2300);
   U227 : AO3 port map( A => n1075, B => n2269, C => n2302, D => n2303, Z => 
                           n6680);
   U228 : AO2 port map( A => n2272, B => v_KEY32_IN_15_port, C => 
                           v_TEMP_VECTOR_23_port, D => n2273, Z => n2303);
   U229 : NR2 port map( A => n2304, B => n2305, Z => n2273);
   U230 : NR2 port map( A => n2305, B => n2306, Z => n2272);
   U231 : MUX21L port map( A => n2307, B => n2308, S => v_TEMP_VECTOR_15_port, 
                           Z => n2302);
   U232 : AO7 port map( A => v_KEY_COL_OUT0_15_port, B => n2276, C => n2277, Z 
                           => n2308);
   U233 : NR2 port map( A => n2276, B => n1068, Z => n2307);
   U234 : OR3 port map( A => n2309, B => n2305, C => n2310, Z => n2276);
   U235 : ND3 port map( A => n2309, B => n2143, C => n2277, Z => n2269);
   U236 : IV port map( A => n2305, Z => n2277);
   U237 : AO7 port map( A => n2311, B => n2309, C => n2156, Z => n2305);
   U238 : AO3 port map( A => n1074, B => n2312, C => n2313, D => n2314, Z => 
                           n6679);
   U239 : AO2 port map( A => n2315, B => v_KEY32_IN_16_port, C => 
                           v_TEMP_VECTOR_24_port, D => n2316, Z => n2314);
   U240 : MUX21L port map( A => n2317, B => n2318, S => v_TEMP_VECTOR_16_port, 
                           Z => n2313);
   U241 : AO7 port map( A => v_KEY_COL_OUT0_16_port, B => n2319, C => n2320, Z 
                           => n2318);
   U242 : NR2 port map( A => n2319, B => n1067, Z => n2317);
   U243 : AO3 port map( A => n4456, B => n2312, C => n2321, D => n2322, Z => 
                           n6678);
   U244 : AO2 port map( A => n2315, B => v_KEY32_IN_17_port, C => 
                           v_TEMP_VECTOR_25_port, D => n2316, Z => n2322);
   U245 : MUX21L port map( A => n2323, B => n2324, S => v_TEMP_VECTOR_17_port, 
                           Z => n2321);
   U246 : AO7 port map( A => v_KEY_COL_OUT0_17_port, B => n2319, C => n2320, Z 
                           => n2324);
   U247 : NR2 port map( A => n2319, B => n1066, Z => n2323);
   U248 : AO3 port map( A => n4465, B => n2312, C => n2325, D => n2326, Z => 
                           n6677);
   U249 : AO2 port map( A => n2315, B => v_KEY32_IN_18_port, C => 
                           v_TEMP_VECTOR_26_port, D => n2316, Z => n2326);
   U250 : MUX21L port map( A => n2327, B => n2328, S => v_TEMP_VECTOR_18_port, 
                           Z => n2325);
   U251 : AO7 port map( A => v_KEY_COL_OUT0_18_port, B => n2319, C => n2320, Z 
                           => n2328);
   U252 : NR2 port map( A => n2319, B => n1065, Z => n2327);
   U253 : AO3 port map( A => n4466, B => n2312, C => n2329, D => n2330, Z => 
                           n6676);
   U254 : AO2 port map( A => n2315, B => v_KEY32_IN_19_port, C => 
                           v_TEMP_VECTOR_27_port, D => n2316, Z => n2330);
   U255 : MUX21L port map( A => n2331, B => n2332, S => v_TEMP_VECTOR_19_port, 
                           Z => n2329);
   U256 : AO7 port map( A => v_KEY_COL_OUT0_19_port, B => n2319, C => n2320, Z 
                           => n2332);
   U257 : NR2 port map( A => n2319, B => n1064, Z => n2331);
   U258 : AO3 port map( A => n4467, B => n2312, C => n2333, D => n2334, Z => 
                           n6675);
   U259 : AO2 port map( A => n2315, B => v_KEY32_IN_20_port, C => 
                           v_TEMP_VECTOR_28_port, D => n2316, Z => n2334);
   U260 : MUX21L port map( A => n2335, B => n2336, S => v_TEMP_VECTOR_20_port, 
                           Z => n2333);
   U261 : AO7 port map( A => v_KEY_COL_OUT0_20_port, B => n2319, C => n2320, Z 
                           => n2336);
   U262 : NR2 port map( A => n2319, B => n1062, Z => n2335);
   U263 : AO3 port map( A => n4468, B => n2312, C => n2337, D => n2338, Z => 
                           n6674);
   U264 : AO2 port map( A => n2315, B => v_KEY32_IN_21_port, C => 
                           v_TEMP_VECTOR_29_port, D => n2316, Z => n2338);
   U265 : MUX21L port map( A => n2339, B => n2340, S => v_TEMP_VECTOR_21_port, 
                           Z => n2337);
   U266 : AO7 port map( A => v_KEY_COL_OUT0_21_port, B => n2319, C => n2320, Z 
                           => n2340);
   U267 : ND2 port map( A => n2319, B => n1061, Z => n2339);
   U268 : AO3 port map( A => n1041, B => n2312, C => n2341, D => n2342, Z => 
                           n6673);
   U269 : AO2 port map( A => n2315, B => v_KEY32_IN_22_port, C => 
                           v_TEMP_VECTOR_30_port, D => n2316, Z => n2342);
   U270 : MUX21L port map( A => n2343, B => n2344, S => v_TEMP_VECTOR_22_port, 
                           Z => n2341);
   U271 : AO7 port map( A => v_KEY_COL_OUT0_22_port, B => n2319, C => n2320, Z 
                           => n2344);
   U272 : ND2 port map( A => n2319, B => n1060, Z => n2343);
   U273 : AO3 port map( A => n1075, B => n2312, C => n2345, D => n2346, Z => 
                           n6672);
   U274 : AO2 port map( A => n2315, B => v_KEY32_IN_23_port, C => 
                           v_TEMP_VECTOR_31_port, D => n2316, Z => n2346);
   U275 : NR2 port map( A => n2347, B => n2304, Z => n2316);
   U276 : NR2 port map( A => n2347, B => n2306, Z => n2315);
   U277 : MUX21L port map( A => n2348, B => n2349, S => v_TEMP_VECTOR_23_port, 
                           Z => n2345);
   U278 : AO7 port map( A => v_KEY_COL_OUT0_23_port, B => n2319, C => n2320, Z 
                           => n2349);
   U279 : NR2 port map( A => n2319, B => n1059, Z => n2348);
   U280 : OR3 port map( A => n2310, B => n2350, C => n2347, Z => n2319);
   U281 : ND3 port map( A => n2350, B => n2143, C => n2320, Z => n2312);
   U282 : IV port map( A => n2347, Z => n2320);
   U283 : AO7 port map( A => n2311, B => n2350, C => n2156, Z => n2347);
   U284 : AO3 port map( A => n1074, B => n2351, C => n2352, D => n2353, Z => 
                           n6671);
   U285 : AO2 port map( A => n2354, B => v_KEY32_IN_24_port, C => n2355, D => 
                           v_TEMP_VECTOR_0_port, Z => n2353);
   U286 : MUX21L port map( A => n2356, B => n2357, S => v_TEMP_VECTOR_24_port, 
                           Z => n2352);
   U287 : AO7 port map( A => v_KEY_COL_OUT0_24_port, B => n2358, C => n2359, Z 
                           => n2357);
   U288 : NR2 port map( A => n2358, B => n1058, Z => n2356);
   U289 : AO3 port map( A => n4456, B => n2351, C => n2360, D => n2361, Z => 
                           n6670);
   U290 : AO2 port map( A => n2354, B => v_KEY32_IN_25_port, C => n2355, D => 
                           v_TEMP_VECTOR_1_port, Z => n2361);
   U291 : MUX21L port map( A => n2362, B => n2363, S => v_TEMP_VECTOR_25_port, 
                           Z => n2360);
   U292 : AO7 port map( A => v_KEY_COL_OUT0_25_port, B => n2358, C => n2359, Z 
                           => n2363);
   U293 : NR2 port map( A => n2358, B => n1057, Z => n2362);
   U294 : AO3 port map( A => n4465, B => n2351, C => n2364, D => n2365, Z => 
                           n6669);
   U295 : AO2 port map( A => n2354, B => v_KEY32_IN_26_port, C => n2355, D => 
                           v_TEMP_VECTOR_2_port, Z => n2365);
   U296 : MUX21L port map( A => n2366, B => n2367, S => v_TEMP_VECTOR_26_port, 
                           Z => n2364);
   U297 : AO7 port map( A => v_KEY_COL_OUT0_26_port, B => n2358, C => n2359, Z 
                           => n2367);
   U298 : NR2 port map( A => n2358, B => n1056, Z => n2366);
   U299 : AO3 port map( A => n4466, B => n2351, C => n2368, D => n2369, Z => 
                           n6668);
   U300 : AO2 port map( A => n2354, B => v_KEY32_IN_27_port, C => n2355, D => 
                           v_TEMP_VECTOR_3_port, Z => n2369);
   U301 : MUX21L port map( A => n2370, B => n2371, S => v_TEMP_VECTOR_27_port, 
                           Z => n2368);
   U302 : AO7 port map( A => v_KEY_COL_OUT0_27_port, B => n2358, C => n2359, Z 
                           => n2371);
   U303 : NR2 port map( A => n2358, B => n1055, Z => n2370);
   U304 : AO3 port map( A => n4467, B => n2351, C => n2372, D => n2373, Z => 
                           n6667);
   U305 : AO2 port map( A => n2354, B => v_KEY32_IN_28_port, C => n2355, D => 
                           v_TEMP_VECTOR_4_port, Z => n2373);
   U306 : MUX21L port map( A => n2374, B => n2375, S => v_TEMP_VECTOR_28_port, 
                           Z => n2372);
   U307 : AO7 port map( A => v_KEY_COL_OUT0_28_port, B => n2358, C => n2359, Z 
                           => n2375);
   U308 : NR2 port map( A => n2358, B => n1054, Z => n2374);
   U309 : AO3 port map( A => n4468, B => n2351, C => n2376, D => n2377, Z => 
                           n6666);
   U310 : AO2 port map( A => n2354, B => v_KEY32_IN_29_port, C => n2355, D => 
                           v_TEMP_VECTOR_5_port, Z => n2377);
   U311 : MUX21L port map( A => n2378, B => n2379, S => v_TEMP_VECTOR_29_port, 
                           Z => n2376);
   U312 : AO7 port map( A => v_KEY_COL_OUT0_29_port, B => n2358, C => n2359, Z 
                           => n2379);
   U313 : NR2 port map( A => n2358, B => n1053, Z => n2378);
   U314 : AO3 port map( A => n1041, B => n2351, C => n2380, D => n2381, Z => 
                           n6665);
   U315 : AO2 port map( A => n2354, B => v_KEY32_IN_30_port, C => n2355, D => 
                           v_TEMP_VECTOR_6_port, Z => n2381);
   U316 : MUX21L port map( A => n2382, B => n2383, S => v_TEMP_VECTOR_30_port, 
                           Z => n2380);
   U317 : AO7 port map( A => v_KEY_COL_OUT0_30_port, B => n2358, C => n2359, Z 
                           => n2383);
   U318 : NR2 port map( A => n2358, B => n1051, Z => n2382);
   U319 : AO3 port map( A => n1075, B => n2351, C => n2384, D => n2385, Z => 
                           n6664);
   U320 : AO2 port map( A => n2354, B => v_KEY32_IN_31_port, C => n2355, D => 
                           v_TEMP_VECTOR_7_port, Z => n2385);
   U321 : NR2 port map( A => n2386, B => n2304, Z => n2355);
   U322 : ND2 port map( A => n2187, B => n2143, Z => n2304);
   U323 : NR2 port map( A => n2386, B => n2306, Z => n2354);
   U324 : IV port map( A => n2266, Z => n2306);
   U325 : NR2 port map( A => n1043, B => RESET_I, Z => n2266);
   U326 : MUX21L port map( A => n2387, B => n2388, S => v_TEMP_VECTOR_31_port, 
                           Z => n2384);
   U327 : AO7 port map( A => v_KEY_COL_OUT0_31_port, B => n2358, C => n2359, Z 
                           => n2388);
   U328 : NR2 port map( A => n2358, B => n1050, Z => n2387);
   U329 : OR3 port map( A => n2310, B => n2389, C => n2386, Z => n2358);
   U330 : ND2 port map( A => n2143, B => n2262, Z => n2310);
   U331 : ND3 port map( A => n2389, B => n2143, C => n2359, Z => n2351);
   U332 : IV port map( A => n2386, Z => n2359);
   U333 : AO7 port map( A => n2311, B => n2389, C => n2156, Z => n2386);
   U334 : ND2 port map( A => n2267, B => n2140, Z => n2156);
   U335 : OR3 port map( A => n2155, B => n2187, C => n2192, Z => n2311);
   U336 : AO4 port map( A => v_CALCULATION_CNTR_2_port, B => n2189, C => n2390,
                           D => n2190, Z => n2192);
   U337 : IV port map( A => n2262, Z => n2187);
   U338 : ND2 port map( A => n2391, B => n2392, Z => n2262);
   U339 : IV port map( A => n2267, Z => n2155);
   U340 : AO6 port map( A => CE_I, B => n4471, C => RESET_I, Z => n2267);
   U341 : IV port map( A => n2153, Z => n2143);
   U342 : MUX21H port map( A => n2393, B => n2394, S => n1036, Z => n2389);
   U343 : NR2 port map( A => n2190, B => n2395, Z => n2394);
   U344 : IV port map( A => n2396, Z => n2190);
   U345 : NR2 port map( A => n2397, B => n2398, Z => n2393);
   U346 : MUX21L port map( A => n2399, B => n2400, S => n8, Z => n6655);
   U347 : ND3 port map( A => v_CALCULATION_CNTR_3_port, B => n2392, C => n2128,
                           Z => n2400);
   U348 : AO6 port map( A => n2128, B => n1078, C => n2401, Z => n2399);
   U349 : IV port map( A => n2402, Z => n2401);
   U350 : MUX21L port map( A => n2403, B => n2402, S => 
                           v_CALCULATION_CNTR_3_port, Z => n6654);
   U351 : AO6 port map( A => n2137, B => n2128, C => n2404, Z => n2402);
   U352 : ND2 port map( A => n2128, B => n2392, Z => n2403);
   U353 : IV port map( A => n2137, Z => n2392);
   U354 : MUX21L port map( A => n2405, B => n2406, S => 
                           v_CALCULATION_CNTR_2_port, Z => n6653);
   U355 : AO6 port map( A => n2128, B => n2407, C => n2404, Z => n2406);
   U356 : ND2 port map( A => n2128, B => n2188, Z => n2405);
   U357 : EON1 port map( A => n7, B => n2136, C => n2408, D => n2128, Z => 
                           n6652);
   U358 : AO7 port map( A => n1077, B => v_CALCULATION_CNTR_1_port, C => n2398,
                           Z => n2408);
   U359 : MUX21L port map( A => n2134, B => n2136, S => 
                           v_CALCULATION_CNTR_0_port, Z => n6651);
   U360 : IV port map( A => n2128, Z => n2134);
   U361 : NR4 port map( A => n2153, B => n2154, C => n2404, D => n4455, Z => 
                           n2128);
   U362 : IV port map( A => n2136, Z => n2404);
   U363 : ND2 port map( A => n2140, B => n2164, Z => n2136);
   U364 : IV port map( A => n2409, Z => n2154);
   U365 : ND2 port map( A => n1043, B => n2164, Z => n2153);
   U366 : IV port map( A => RESET_I, Z => n2164);
   U367 : MUX21L port map( A => n2410, B => n1131, S => n2411, Z => n6637);
   U368 : MUX21L port map( A => n2410, B => n60, S => n2412, Z => n6636);
   U369 : MUX21L port map( A => n2410, B => n1130, S => n2413, Z => n6635);
   U370 : MUX21L port map( A => n2410, B => n59, S => n2414, Z => n6634);
   U371 : MUX21L port map( A => n1129, B => n2410, S => n2415, Z => n6633);
   U372 : MUX21L port map( A => n58, B => n2410, S => n2416, Z => n6632);
   U373 : MUX21L port map( A => n1128, B => n2410, S => n2417, Z => n6631);
   U374 : MUX21L port map( A => n57, B => n2410, S => n2418, Z => n6630);
   U375 : MUX21L port map( A => n2410, B => n1135, S => n2419, Z => n6629);
   U376 : MUX21L port map( A => n2410, B => n64, S => n2420, Z => n6628);
   U377 : MUX21L port map( A => n2410, B => n1134, S => n2421, Z => n6627);
   U378 : MUX21L port map( A => n2410, B => n63, S => n2422, Z => n6626);
   U379 : MUX21L port map( A => n1133, B => n2410, S => n2423, Z => n6625);
   U380 : MUX21L port map( A => n62, B => n2410, S => n2424, Z => n6624);
   U381 : MUX21L port map( A => n1132, B => n2410, S => n2425, Z => n6623);
   U382 : MUX21L port map( A => n61, B => n2410, S => n2426, Z => n6622);
   U383 : MUX21L port map( A => n2410, B => n1139, S => n2427, Z => n6621);
   U384 : MUX21L port map( A => n2410, B => n68, S => n2428, Z => n6620);
   U385 : MUX21L port map( A => n2410, B => n1138, S => n2429, Z => n6619);
   U386 : MUX21L port map( A => n2410, B => n67, S => n2430, Z => n6618);
   U387 : MUX21L port map( A => n1137, B => n2410, S => n2431, Z => n6617);
   U388 : MUX21L port map( A => n66, B => n2410, S => n2432, Z => n6616);
   U389 : MUX21L port map( A => n1136, B => n2410, S => n2433, Z => n6615);
   U390 : MUX21L port map( A => n65, B => n2410, S => n2434, Z => n6614);
   U391 : MUX21L port map( A => n2410, B => n1143, S => n2435, Z => n6613);
   U392 : MUX21L port map( A => n2410, B => n72, S => n2436, Z => n6612);
   U393 : MUX21L port map( A => n2410, B => n1142, S => n2437, Z => n6611);
   U394 : MUX21L port map( A => n2410, B => n71, S => n2438, Z => n6610);
   U395 : MUX21L port map( A => n1141, B => n2410, S => n2439, Z => n6609);
   U396 : MUX21L port map( A => n70, B => n2410, S => n2440, Z => n6608);
   U397 : MUX21L port map( A => n1140, B => n2410, S => n2441, Z => n6607);
   U398 : MUX21L port map( A => n69, B => n2410, S => n2442, Z => n6606);
   U399 : MUX21L port map( A => n2410, B => n1115, S => n2443, Z => n6605);
   U400 : MUX21L port map( A => n2410, B => n44, S => n2444, Z => n6604);
   U401 : MUX21L port map( A => n2410, B => n1114, S => n2445, Z => n6603);
   U402 : MUX21L port map( A => n2410, B => n43, S => n2446, Z => n6602);
   U403 : MUX21L port map( A => n1113, B => n2410, S => n2447, Z => n6601);
   U404 : MUX21L port map( A => n42, B => n2410, S => n2448, Z => n6600);
   U405 : MUX21L port map( A => n1112, B => n2410, S => n2449, Z => n6599);
   U406 : MUX21L port map( A => n41, B => n2410, S => n2450, Z => n6598);
   U407 : MUX21L port map( A => n2410, B => n1119, S => n2451, Z => n6597);
   U408 : MUX21L port map( A => n2410, B => n48, S => n2452, Z => n6596);
   U409 : MUX21L port map( A => n2410, B => n1118, S => n2453, Z => n6595);
   U410 : MUX21L port map( A => n2410, B => n47, S => n2454, Z => n6594);
   U411 : MUX21L port map( A => n1117, B => n2410, S => n2455, Z => n6593);
   U412 : MUX21L port map( A => n46, B => n2410, S => n2456, Z => n6592);
   U413 : MUX21L port map( A => n1116, B => n2410, S => n2457, Z => n6591);
   U414 : MUX21L port map( A => n45, B => n2410, S => n2458, Z => n6590);
   U415 : MUX21L port map( A => n2410, B => n1123, S => n2459, Z => n6589);
   U416 : MUX21L port map( A => n2410, B => n52, S => n2460, Z => n6588);
   U417 : MUX21L port map( A => n2410, B => n1122, S => n2461, Z => n6587);
   U418 : MUX21L port map( A => n2410, B => n51, S => n2462, Z => n6586);
   U419 : MUX21L port map( A => n1121, B => n2410, S => n2463, Z => n6585);
   U420 : MUX21L port map( A => n50, B => n2410, S => n2464, Z => n6584);
   U421 : MUX21L port map( A => n1120, B => n2410, S => n2465, Z => n6583);
   U422 : MUX21L port map( A => n49, B => n2410, S => n2466, Z => n6582);
   U423 : MUX21L port map( A => n2410, B => n1127, S => n2467, Z => n6581);
   U424 : MUX21L port map( A => n2410, B => n56, S => n2468, Z => n6580);
   U425 : MUX21L port map( A => n2410, B => n1126, S => n2469, Z => n6579);
   U426 : MUX21L port map( A => n2410, B => n55, S => n2470, Z => n6578);
   U427 : MUX21L port map( A => n1125, B => n2410, S => n2471, Z => n6577);
   U428 : MUX21L port map( A => n54, B => n2410, S => n2472, Z => n6576);
   U429 : MUX21L port map( A => n1124, B => n2410, S => n2473, Z => n6575);
   U430 : MUX21L port map( A => n53, B => n2410, S => n2474, Z => n6574);
   U431 : AO2 port map( A => v_TEMP_VECTOR_31_port, B => n2475, C => 
                           v_KEY32_IN_31_port, D => n2476, Z => n2410);
   U432 : MUX21L port map( A => n2477, B => n1259, S => n2411, Z => n6573);
   U433 : MUX21L port map( A => n2477, B => n188, S => n2412, Z => n6572);
   U434 : MUX21L port map( A => n2477, B => n1258, S => n2413, Z => n6571);
   U435 : MUX21L port map( A => n2477, B => n187, S => n2414, Z => n6570);
   U436 : MUX21L port map( A => n1257, B => n2477, S => n2415, Z => n6569);
   U437 : MUX21L port map( A => n186, B => n2477, S => n2416, Z => n6568);
   U438 : MUX21L port map( A => n1256, B => n2477, S => n2417, Z => n6567);
   U439 : MUX21L port map( A => n185, B => n2477, S => n2418, Z => n6566);
   U440 : MUX21L port map( A => n2477, B => n1263, S => n2419, Z => n6565);
   U441 : MUX21L port map( A => n2477, B => n192, S => n2420, Z => n6564);
   U442 : MUX21L port map( A => n2477, B => n1262, S => n2421, Z => n6563);
   U443 : MUX21L port map( A => n2477, B => n191, S => n2422, Z => n6562);
   U444 : MUX21L port map( A => n1261, B => n2477, S => n2423, Z => n6561);
   U445 : MUX21L port map( A => n190, B => n2477, S => n2424, Z => n6560);
   U446 : MUX21L port map( A => n1260, B => n2477, S => n2425, Z => n6559);
   U447 : MUX21L port map( A => n189, B => n2477, S => n2426, Z => n6558);
   U448 : MUX21L port map( A => n2477, B => n1267, S => n2427, Z => n6557);
   U449 : MUX21L port map( A => n2477, B => n196, S => n2428, Z => n6556);
   U450 : MUX21L port map( A => n2477, B => n1266, S => n2429, Z => n6555);
   U451 : MUX21L port map( A => n2477, B => n195, S => n2430, Z => n6554);
   U452 : MUX21L port map( A => n1265, B => n2477, S => n2431, Z => n6553);
   U453 : MUX21L port map( A => n194, B => n2477, S => n2432, Z => n6552);
   U454 : MUX21L port map( A => n1264, B => n2477, S => n2433, Z => n6551);
   U455 : MUX21L port map( A => n193, B => n2477, S => n2434, Z => n6550);
   U456 : MUX21L port map( A => n2477, B => n1271, S => n2435, Z => n6549);
   U457 : MUX21L port map( A => n2477, B => n200, S => n2436, Z => n6548);
   U458 : MUX21L port map( A => n2477, B => n1270, S => n2437, Z => n6547);
   U459 : MUX21L port map( A => n2477, B => n199, S => n2438, Z => n6546);
   U460 : MUX21L port map( A => n1269, B => n2477, S => n2439, Z => n6545);
   U461 : MUX21L port map( A => n198, B => n2477, S => n2440, Z => n6544);
   U462 : MUX21L port map( A => n1268, B => n2477, S => n2441, Z => n6543);
   U463 : MUX21L port map( A => n197, B => n2477, S => n2442, Z => n6542);
   U464 : MUX21L port map( A => n2477, B => n1243, S => n2443, Z => n6541);
   U465 : MUX21L port map( A => n2477, B => n172, S => n2444, Z => n6540);
   U466 : MUX21L port map( A => n2477, B => n1242, S => n2445, Z => n6539);
   U467 : MUX21L port map( A => n2477, B => n171, S => n2446, Z => n6538);
   U468 : MUX21L port map( A => n1241, B => n2477, S => n2447, Z => n6537);
   U469 : MUX21L port map( A => n170, B => n2477, S => n2448, Z => n6536);
   U470 : MUX21L port map( A => n1240, B => n2477, S => n2449, Z => n6535);
   U471 : MUX21L port map( A => n169, B => n2477, S => n2450, Z => n6534);
   U472 : MUX21L port map( A => n2477, B => n1247, S => n2451, Z => n6533);
   U473 : MUX21L port map( A => n2477, B => n176, S => n2452, Z => n6532);
   U474 : MUX21L port map( A => n2477, B => n1246, S => n2453, Z => n6531);
   U475 : MUX21L port map( A => n2477, B => n175, S => n2454, Z => n6530);
   U476 : MUX21L port map( A => n1245, B => n2477, S => n2455, Z => n6529);
   U477 : MUX21L port map( A => n174, B => n2477, S => n2456, Z => n6528);
   U478 : MUX21L port map( A => n1244, B => n2477, S => n2457, Z => n6527);
   U479 : MUX21L port map( A => n173, B => n2477, S => n2458, Z => n6526);
   U480 : MUX21L port map( A => n2477, B => n1251, S => n2459, Z => n6525);
   U481 : MUX21L port map( A => n2477, B => n180, S => n2460, Z => n6524);
   U482 : MUX21L port map( A => n2477, B => n1250, S => n2461, Z => n6523);
   U483 : MUX21L port map( A => n2477, B => n179, S => n2462, Z => n6522);
   U484 : MUX21L port map( A => n1249, B => n2477, S => n2463, Z => n6521);
   U485 : MUX21L port map( A => n178, B => n2477, S => n2464, Z => n6520);
   U486 : MUX21L port map( A => n1248, B => n2477, S => n2465, Z => n6519);
   U487 : MUX21L port map( A => n177, B => n2477, S => n2466, Z => n6518);
   U488 : MUX21L port map( A => n2477, B => n1255, S => n2467, Z => n6517);
   U489 : MUX21L port map( A => n2477, B => n184, S => n2468, Z => n6516);
   U490 : MUX21L port map( A => n2477, B => n1254, S => n2469, Z => n6515);
   U491 : MUX21L port map( A => n2477, B => n183, S => n2470, Z => n6514);
   U492 : MUX21L port map( A => n1253, B => n2477, S => n2471, Z => n6513);
   U493 : MUX21L port map( A => n182, B => n2477, S => n2472, Z => n6512);
   U494 : MUX21L port map( A => n1252, B => n2477, S => n2473, Z => n6511);
   U495 : MUX21L port map( A => n181, B => n2477, S => n2474, Z => n6510);
   U496 : AO2 port map( A => v_TEMP_VECTOR_30_port, B => n2475, C => 
                           v_KEY32_IN_30_port, D => n2476, Z => n2477);
   U497 : MUX21L port map( A => n2478, B => n1387, S => n2411, Z => n6509);
   U498 : MUX21L port map( A => n2478, B => n316, S => n2412, Z => n6508);
   U499 : MUX21L port map( A => n2478, B => n1386, S => n2413, Z => n6507);
   U500 : MUX21L port map( A => n2478, B => n315, S => n2414, Z => n6506);
   U501 : MUX21L port map( A => n1385, B => n2478, S => n2415, Z => n6505);
   U502 : MUX21L port map( A => n314, B => n2478, S => n2416, Z => n6504);
   U503 : MUX21L port map( A => n1384, B => n2478, S => n2417, Z => n6503);
   U504 : MUX21L port map( A => n313, B => n2478, S => n2418, Z => n6502);
   U505 : MUX21L port map( A => n2478, B => n1391, S => n2419, Z => n6501);
   U506 : MUX21L port map( A => n2478, B => n320, S => n2420, Z => n6500);
   U507 : MUX21L port map( A => n2478, B => n1390, S => n2421, Z => n6499);
   U508 : MUX21L port map( A => n2478, B => n319, S => n2422, Z => n6498);
   U509 : MUX21L port map( A => n1389, B => n2478, S => n2423, Z => n6497);
   U510 : MUX21L port map( A => n318, B => n2478, S => n2424, Z => n6496);
   U511 : MUX21L port map( A => n1388, B => n2478, S => n2425, Z => n6495);
   U512 : MUX21L port map( A => n317, B => n2478, S => n2426, Z => n6494);
   U513 : MUX21L port map( A => n2478, B => n1395, S => n2427, Z => n6493);
   U514 : MUX21L port map( A => n2478, B => n324, S => n2428, Z => n6492);
   U515 : MUX21L port map( A => n2478, B => n1394, S => n2429, Z => n6491);
   U516 : MUX21L port map( A => n2478, B => n323, S => n2430, Z => n6490);
   U517 : MUX21L port map( A => n1393, B => n2478, S => n2431, Z => n6489);
   U518 : MUX21L port map( A => n322, B => n2478, S => n2432, Z => n6488);
   U519 : MUX21L port map( A => n1392, B => n2478, S => n2433, Z => n6487);
   U520 : MUX21L port map( A => n321, B => n2478, S => n2434, Z => n6486);
   U521 : MUX21L port map( A => n2478, B => n1399, S => n2435, Z => n6485);
   U522 : MUX21L port map( A => n2478, B => n328, S => n2436, Z => n6484);
   U523 : MUX21L port map( A => n2478, B => n1398, S => n2437, Z => n6483);
   U524 : MUX21L port map( A => n2478, B => n327, S => n2438, Z => n6482);
   U525 : MUX21L port map( A => n1397, B => n2478, S => n2439, Z => n6481);
   U526 : MUX21L port map( A => n326, B => n2478, S => n2440, Z => n6480);
   U527 : MUX21L port map( A => n1396, B => n2478, S => n2441, Z => n6479);
   U528 : MUX21L port map( A => n325, B => n2478, S => n2442, Z => n6478);
   U529 : MUX21L port map( A => n2478, B => n1371, S => n2443, Z => n6477);
   U530 : MUX21L port map( A => n2478, B => n300, S => n2444, Z => n6476);
   U531 : MUX21L port map( A => n2478, B => n1370, S => n2445, Z => n6475);
   U532 : MUX21L port map( A => n2478, B => n299, S => n2446, Z => n6474);
   U533 : MUX21L port map( A => n1369, B => n2478, S => n2447, Z => n6473);
   U534 : MUX21L port map( A => n298, B => n2478, S => n2448, Z => n6472);
   U535 : MUX21L port map( A => n1368, B => n2478, S => n2449, Z => n6471);
   U536 : MUX21L port map( A => n297, B => n2478, S => n2450, Z => n6470);
   U537 : MUX21L port map( A => n2478, B => n1375, S => n2451, Z => n6469);
   U538 : MUX21L port map( A => n2478, B => n304, S => n2452, Z => n6468);
   U539 : MUX21L port map( A => n2478, B => n1374, S => n2453, Z => n6467);
   U540 : MUX21L port map( A => n2478, B => n303, S => n2454, Z => n6466);
   U541 : MUX21L port map( A => n1373, B => n2478, S => n2455, Z => n6465);
   U542 : MUX21L port map( A => n302, B => n2478, S => n2456, Z => n6464);
   U543 : MUX21L port map( A => n1372, B => n2478, S => n2457, Z => n6463);
   U544 : MUX21L port map( A => n301, B => n2478, S => n2458, Z => n6462);
   U545 : MUX21L port map( A => n2478, B => n1379, S => n2459, Z => n6461);
   U546 : MUX21L port map( A => n2478, B => n308, S => n2460, Z => n6460);
   U547 : MUX21L port map( A => n2478, B => n1378, S => n2461, Z => n6459);
   U548 : MUX21L port map( A => n2478, B => n307, S => n2462, Z => n6458);
   U549 : MUX21L port map( A => n1377, B => n2478, S => n2463, Z => n6457);
   U550 : MUX21L port map( A => n306, B => n2478, S => n2464, Z => n6456);
   U551 : MUX21L port map( A => n1376, B => n2478, S => n2465, Z => n6455);
   U552 : MUX21L port map( A => n305, B => n2478, S => n2466, Z => n6454);
   U553 : MUX21L port map( A => n2478, B => n1383, S => n2467, Z => n6453);
   U554 : MUX21L port map( A => n2478, B => n312, S => n2468, Z => n6452);
   U555 : MUX21L port map( A => n2478, B => n1382, S => n2469, Z => n6451);
   U556 : MUX21L port map( A => n2478, B => n311, S => n2470, Z => n6450);
   U557 : MUX21L port map( A => n1381, B => n2478, S => n2471, Z => n6449);
   U558 : MUX21L port map( A => n310, B => n2478, S => n2472, Z => n6448);
   U559 : MUX21L port map( A => n1380, B => n2478, S => n2473, Z => n6447);
   U560 : MUX21L port map( A => n309, B => n2478, S => n2474, Z => n6446);
   U561 : AO2 port map( A => v_TEMP_VECTOR_29_port, B => n2475, C => 
                           v_KEY32_IN_29_port, D => n2476, Z => n2478);
   U562 : MUX21L port map( A => n2479, B => n1515, S => n2411, Z => n6445);
   U563 : MUX21L port map( A => n2479, B => n444, S => n2412, Z => n6444);
   U564 : MUX21L port map( A => n2479, B => n1514, S => n2413, Z => n6443);
   U565 : MUX21L port map( A => n2479, B => n443, S => n2414, Z => n6442);
   U566 : MUX21L port map( A => n1513, B => n2479, S => n2415, Z => n6441);
   U567 : MUX21L port map( A => n442, B => n2479, S => n2416, Z => n6440);
   U568 : MUX21L port map( A => n1512, B => n2479, S => n2417, Z => n6439);
   U569 : MUX21L port map( A => n441, B => n2479, S => n2418, Z => n6438);
   U570 : MUX21L port map( A => n2479, B => n1519, S => n2419, Z => n6437);
   U571 : MUX21L port map( A => n2479, B => n448, S => n2420, Z => n6436);
   U572 : MUX21L port map( A => n2479, B => n1518, S => n2421, Z => n6435);
   U573 : MUX21L port map( A => n2479, B => n447, S => n2422, Z => n6434);
   U574 : MUX21L port map( A => n1517, B => n2479, S => n2423, Z => n6433);
   U575 : MUX21L port map( A => n446, B => n2479, S => n2424, Z => n6432);
   U576 : MUX21L port map( A => n1516, B => n2479, S => n2425, Z => n6431);
   U577 : MUX21L port map( A => n445, B => n2479, S => n2426, Z => n6430);
   U578 : MUX21L port map( A => n2479, B => n1523, S => n2427, Z => n6429);
   U579 : MUX21L port map( A => n2479, B => n452, S => n2428, Z => n6428);
   U580 : MUX21L port map( A => n2479, B => n1522, S => n2429, Z => n6427);
   U581 : MUX21L port map( A => n2479, B => n451, S => n2430, Z => n6426);
   U582 : MUX21L port map( A => n1521, B => n2479, S => n2431, Z => n6425);
   U583 : MUX21L port map( A => n450, B => n2479, S => n2432, Z => n6424);
   U584 : MUX21L port map( A => n1520, B => n2479, S => n2433, Z => n6423);
   U585 : MUX21L port map( A => n449, B => n2479, S => n2434, Z => n6422);
   U586 : MUX21L port map( A => n2479, B => n1527, S => n2435, Z => n6421);
   U587 : MUX21L port map( A => n2479, B => n456, S => n2436, Z => n6420);
   U588 : MUX21L port map( A => n2479, B => n1526, S => n2437, Z => n6419);
   U589 : MUX21L port map( A => n2479, B => n455, S => n2438, Z => n6418);
   U590 : MUX21L port map( A => n1525, B => n2479, S => n2439, Z => n6417);
   U591 : MUX21L port map( A => n454, B => n2479, S => n2440, Z => n6416);
   U592 : MUX21L port map( A => n1524, B => n2479, S => n2441, Z => n6415);
   U593 : MUX21L port map( A => n453, B => n2479, S => n2442, Z => n6414);
   U594 : MUX21L port map( A => n2479, B => n1499, S => n2443, Z => n6413);
   U595 : MUX21L port map( A => n2479, B => n428, S => n2444, Z => n6412);
   U596 : MUX21L port map( A => n2479, B => n1498, S => n2445, Z => n6411);
   U597 : MUX21L port map( A => n2479, B => n427, S => n2446, Z => n6410);
   U598 : MUX21L port map( A => n1497, B => n2479, S => n2447, Z => n6409);
   U599 : MUX21L port map( A => n426, B => n2479, S => n2448, Z => n6408);
   U600 : MUX21L port map( A => n1496, B => n2479, S => n2449, Z => n6407);
   U601 : MUX21L port map( A => n425, B => n2479, S => n2450, Z => n6406);
   U602 : MUX21L port map( A => n2479, B => n1503, S => n2451, Z => n6405);
   U603 : MUX21L port map( A => n2479, B => n432, S => n2452, Z => n6404);
   U604 : MUX21L port map( A => n2479, B => n1502, S => n2453, Z => n6403);
   U605 : MUX21L port map( A => n2479, B => n431, S => n2454, Z => n6402);
   U606 : MUX21L port map( A => n1501, B => n2479, S => n2455, Z => n6401);
   U607 : MUX21L port map( A => n430, B => n2479, S => n2456, Z => n6400);
   U608 : MUX21L port map( A => n1500, B => n2479, S => n2457, Z => n6399);
   U609 : MUX21L port map( A => n429, B => n2479, S => n2458, Z => n6398);
   U610 : MUX21L port map( A => n2479, B => n1507, S => n2459, Z => n6397);
   U611 : MUX21L port map( A => n2479, B => n436, S => n2460, Z => n6396);
   U612 : MUX21L port map( A => n2479, B => n1506, S => n2461, Z => n6395);
   U613 : MUX21L port map( A => n2479, B => n435, S => n2462, Z => n6394);
   U614 : MUX21L port map( A => n1505, B => n2479, S => n2463, Z => n6393);
   U615 : MUX21L port map( A => n434, B => n2479, S => n2464, Z => n6392);
   U616 : MUX21L port map( A => n1504, B => n2479, S => n2465, Z => n6391);
   U617 : MUX21L port map( A => n433, B => n2479, S => n2466, Z => n6390);
   U618 : MUX21L port map( A => n2479, B => n1511, S => n2467, Z => n6389);
   U619 : MUX21L port map( A => n2479, B => n440, S => n2468, Z => n6388);
   U620 : MUX21L port map( A => n2479, B => n1510, S => n2469, Z => n6387);
   U621 : MUX21L port map( A => n2479, B => n439, S => n2470, Z => n6386);
   U622 : MUX21L port map( A => n1509, B => n2479, S => n2471, Z => n6385);
   U623 : MUX21L port map( A => n438, B => n2479, S => n2472, Z => n6384);
   U624 : MUX21L port map( A => n1508, B => n2479, S => n2473, Z => n6383);
   U625 : MUX21L port map( A => n437, B => n2479, S => n2474, Z => n6382);
   U626 : AO2 port map( A => v_TEMP_VECTOR_28_port, B => n2475, C => 
                           v_KEY32_IN_28_port, D => n2476, Z => n2479);
   U627 : MUX21L port map( A => n2480, B => n1643, S => n2411, Z => n6381);
   U628 : MUX21L port map( A => n2480, B => n572, S => n2412, Z => n6380);
   U629 : MUX21L port map( A => n2480, B => n1642, S => n2413, Z => n6379);
   U630 : MUX21L port map( A => n2480, B => n571, S => n2414, Z => n6378);
   U631 : MUX21L port map( A => n1641, B => n2480, S => n2415, Z => n6377);
   U632 : MUX21L port map( A => n570, B => n2480, S => n2416, Z => n6376);
   U633 : MUX21L port map( A => n1640, B => n2480, S => n2417, Z => n6375);
   U634 : MUX21L port map( A => n569, B => n2480, S => n2418, Z => n6374);
   U635 : MUX21L port map( A => n2480, B => n1647, S => n2419, Z => n6373);
   U636 : MUX21L port map( A => n2480, B => n576, S => n2420, Z => n6372);
   U637 : MUX21L port map( A => n2480, B => n1646, S => n2421, Z => n6371);
   U638 : MUX21L port map( A => n2480, B => n575, S => n2422, Z => n6370);
   U639 : MUX21L port map( A => n1645, B => n2480, S => n2423, Z => n6369);
   U640 : MUX21L port map( A => n574, B => n2480, S => n2424, Z => n6368);
   U641 : MUX21L port map( A => n1644, B => n2480, S => n2425, Z => n6367);
   U642 : MUX21L port map( A => n573, B => n2480, S => n2426, Z => n6366);
   U643 : MUX21L port map( A => n2480, B => n1651, S => n2427, Z => n6365);
   U644 : MUX21L port map( A => n2480, B => n580, S => n2428, Z => n6364);
   U645 : MUX21L port map( A => n2480, B => n1650, S => n2429, Z => n6363);
   U646 : MUX21L port map( A => n2480, B => n579, S => n2430, Z => n6362);
   U647 : MUX21L port map( A => n1649, B => n2480, S => n2431, Z => n6361);
   U648 : MUX21L port map( A => n578, B => n2480, S => n2432, Z => n6360);
   U649 : MUX21L port map( A => n1648, B => n2480, S => n2433, Z => n6359);
   U650 : MUX21L port map( A => n577, B => n2480, S => n2434, Z => n6358);
   U651 : MUX21L port map( A => n2480, B => n1655, S => n2435, Z => n6357);
   U652 : MUX21L port map( A => n2480, B => n584, S => n2436, Z => n6356);
   U653 : MUX21L port map( A => n2480, B => n1654, S => n2437, Z => n6355);
   U654 : MUX21L port map( A => n2480, B => n583, S => n2438, Z => n6354);
   U655 : MUX21L port map( A => n1653, B => n2480, S => n2439, Z => n6353);
   U656 : MUX21L port map( A => n582, B => n2480, S => n2440, Z => n6352);
   U657 : MUX21L port map( A => n1652, B => n2480, S => n2441, Z => n6351);
   U658 : MUX21L port map( A => n581, B => n2480, S => n2442, Z => n6350);
   U659 : MUX21L port map( A => n2480, B => n1627, S => n2443, Z => n6349);
   U660 : MUX21L port map( A => n2480, B => n556, S => n2444, Z => n6348);
   U661 : MUX21L port map( A => n2480, B => n1626, S => n2445, Z => n6347);
   U662 : MUX21L port map( A => n2480, B => n555, S => n2446, Z => n6346);
   U663 : MUX21L port map( A => n1625, B => n2480, S => n2447, Z => n6345);
   U664 : MUX21L port map( A => n554, B => n2480, S => n2448, Z => n6344);
   U665 : MUX21L port map( A => n1624, B => n2480, S => n2449, Z => n6343);
   U666 : MUX21L port map( A => n553, B => n2480, S => n2450, Z => n6342);
   U667 : MUX21L port map( A => n2480, B => n1631, S => n2451, Z => n6341);
   U668 : MUX21L port map( A => n2480, B => n560, S => n2452, Z => n6340);
   U669 : MUX21L port map( A => n2480, B => n1630, S => n2453, Z => n6339);
   U670 : MUX21L port map( A => n2480, B => n559, S => n2454, Z => n6338);
   U671 : MUX21L port map( A => n1629, B => n2480, S => n2455, Z => n6337);
   U672 : MUX21L port map( A => n558, B => n2480, S => n2456, Z => n6336);
   U673 : MUX21L port map( A => n1628, B => n2480, S => n2457, Z => n6335);
   U674 : MUX21L port map( A => n557, B => n2480, S => n2458, Z => n6334);
   U675 : MUX21L port map( A => n2480, B => n1635, S => n2459, Z => n6333);
   U676 : MUX21L port map( A => n2480, B => n564, S => n2460, Z => n6332);
   U677 : MUX21L port map( A => n2480, B => n1634, S => n2461, Z => n6331);
   U678 : MUX21L port map( A => n2480, B => n563, S => n2462, Z => n6330);
   U679 : MUX21L port map( A => n1633, B => n2480, S => n2463, Z => n6329);
   U680 : MUX21L port map( A => n562, B => n2480, S => n2464, Z => n6328);
   U681 : MUX21L port map( A => n1632, B => n2480, S => n2465, Z => n6327);
   U682 : MUX21L port map( A => n561, B => n2480, S => n2466, Z => n6326);
   U683 : MUX21L port map( A => n2480, B => n1639, S => n2467, Z => n6325);
   U684 : MUX21L port map( A => n2480, B => n568, S => n2468, Z => n6324);
   U685 : MUX21L port map( A => n2480, B => n1638, S => n2469, Z => n6323);
   U686 : MUX21L port map( A => n2480, B => n567, S => n2470, Z => n6322);
   U687 : MUX21L port map( A => n1637, B => n2480, S => n2471, Z => n6321);
   U688 : MUX21L port map( A => n566, B => n2480, S => n2472, Z => n6320);
   U689 : MUX21L port map( A => n1636, B => n2480, S => n2473, Z => n6319);
   U690 : MUX21L port map( A => n565, B => n2480, S => n2474, Z => n6318);
   U691 : AO2 port map( A => v_TEMP_VECTOR_27_port, B => n2475, C => 
                           v_KEY32_IN_27_port, D => n2476, Z => n2480);
   U692 : MUX21L port map( A => n2481, B => n1771, S => n2411, Z => n6317);
   U693 : MUX21L port map( A => n2481, B => n700, S => n2412, Z => n6316);
   U694 : MUX21L port map( A => n2481, B => n1770, S => n2413, Z => n6315);
   U695 : MUX21L port map( A => n2481, B => n699, S => n2414, Z => n6314);
   U696 : MUX21L port map( A => n1769, B => n2481, S => n2415, Z => n6313);
   U697 : MUX21L port map( A => n698, B => n2481, S => n2416, Z => n6312);
   U698 : MUX21L port map( A => n1768, B => n2481, S => n2417, Z => n6311);
   U699 : MUX21L port map( A => n697, B => n2481, S => n2418, Z => n6310);
   U700 : MUX21L port map( A => n2481, B => n1775, S => n2419, Z => n6309);
   U701 : MUX21L port map( A => n2481, B => n704, S => n2420, Z => n6308);
   U702 : MUX21L port map( A => n2481, B => n1774, S => n2421, Z => n6307);
   U703 : MUX21L port map( A => n2481, B => n703, S => n2422, Z => n6306);
   U704 : MUX21L port map( A => n1773, B => n2481, S => n2423, Z => n6305);
   U705 : MUX21L port map( A => n702, B => n2481, S => n2424, Z => n6304);
   U706 : MUX21L port map( A => n1772, B => n2481, S => n2425, Z => n6303);
   U707 : MUX21L port map( A => n701, B => n2481, S => n2426, Z => n6302);
   U708 : MUX21L port map( A => n2481, B => n1779, S => n2427, Z => n6301);
   U709 : MUX21L port map( A => n2481, B => n708, S => n2428, Z => n6300);
   U710 : MUX21L port map( A => n2481, B => n1778, S => n2429, Z => n6299);
   U711 : MUX21L port map( A => n2481, B => n707, S => n2430, Z => n6298);
   U712 : MUX21L port map( A => n1777, B => n2481, S => n2431, Z => n6297);
   U713 : MUX21L port map( A => n706, B => n2481, S => n2432, Z => n6296);
   U714 : MUX21L port map( A => n1776, B => n2481, S => n2433, Z => n6295);
   U715 : MUX21L port map( A => n705, B => n2481, S => n2434, Z => n6294);
   U716 : MUX21L port map( A => n2481, B => n1783, S => n2435, Z => n6293);
   U717 : MUX21L port map( A => n2481, B => n712, S => n2436, Z => n6292);
   U718 : MUX21L port map( A => n2481, B => n1782, S => n2437, Z => n6291);
   U719 : MUX21L port map( A => n2481, B => n711, S => n2438, Z => n6290);
   U720 : MUX21L port map( A => n1781, B => n2481, S => n2439, Z => n6289);
   U721 : MUX21L port map( A => n710, B => n2481, S => n2440, Z => n6288);
   U722 : MUX21L port map( A => n1780, B => n2481, S => n2441, Z => n6287);
   U723 : MUX21L port map( A => n709, B => n2481, S => n2442, Z => n6286);
   U724 : MUX21L port map( A => n2481, B => n1755, S => n2443, Z => n6285);
   U725 : MUX21L port map( A => n2481, B => n684, S => n2444, Z => n6284);
   U726 : MUX21L port map( A => n2481, B => n1754, S => n2445, Z => n6283);
   U727 : MUX21L port map( A => n2481, B => n683, S => n2446, Z => n6282);
   U728 : MUX21L port map( A => n1753, B => n2481, S => n2447, Z => n6281);
   U729 : MUX21L port map( A => n682, B => n2481, S => n2448, Z => n6280);
   U730 : MUX21L port map( A => n1752, B => n2481, S => n2449, Z => n6279);
   U731 : MUX21L port map( A => n681, B => n2481, S => n2450, Z => n6278);
   U732 : MUX21L port map( A => n2481, B => n1759, S => n2451, Z => n6277);
   U733 : MUX21L port map( A => n2481, B => n688, S => n2452, Z => n6276);
   U734 : MUX21L port map( A => n2481, B => n1758, S => n2453, Z => n6275);
   U735 : MUX21L port map( A => n2481, B => n687, S => n2454, Z => n6274);
   U736 : MUX21L port map( A => n1757, B => n2481, S => n2455, Z => n6273);
   U737 : MUX21L port map( A => n686, B => n2481, S => n2456, Z => n6272);
   U738 : MUX21L port map( A => n1756, B => n2481, S => n2457, Z => n6271);
   U739 : MUX21L port map( A => n685, B => n2481, S => n2458, Z => n6270);
   U740 : MUX21L port map( A => n2481, B => n1763, S => n2459, Z => n6269);
   U741 : MUX21L port map( A => n2481, B => n692, S => n2460, Z => n6268);
   U742 : MUX21L port map( A => n2481, B => n1762, S => n2461, Z => n6267);
   U743 : MUX21L port map( A => n2481, B => n691, S => n2462, Z => n6266);
   U744 : MUX21L port map( A => n1761, B => n2481, S => n2463, Z => n6265);
   U745 : MUX21L port map( A => n690, B => n2481, S => n2464, Z => n6264);
   U746 : MUX21L port map( A => n1760, B => n2481, S => n2465, Z => n6263);
   U747 : MUX21L port map( A => n689, B => n2481, S => n2466, Z => n6262);
   U748 : MUX21L port map( A => n2481, B => n1767, S => n2467, Z => n6261);
   U749 : MUX21L port map( A => n2481, B => n696, S => n2468, Z => n6260);
   U750 : MUX21L port map( A => n2481, B => n1766, S => n2469, Z => n6259);
   U751 : MUX21L port map( A => n2481, B => n695, S => n2470, Z => n6258);
   U752 : MUX21L port map( A => n1765, B => n2481, S => n2471, Z => n6257);
   U753 : MUX21L port map( A => n694, B => n2481, S => n2472, Z => n6256);
   U754 : MUX21L port map( A => n1764, B => n2481, S => n2473, Z => n6255);
   U755 : MUX21L port map( A => n693, B => n2481, S => n2474, Z => n6254);
   U756 : AO2 port map( A => v_TEMP_VECTOR_26_port, B => n2475, C => 
                           v_KEY32_IN_26_port, D => n2476, Z => n2481);
   U757 : MUX21L port map( A => n2482, B => n1899, S => n2411, Z => n6253);
   U758 : MUX21L port map( A => n2482, B => n828, S => n2412, Z => n6252);
   U759 : MUX21L port map( A => n2482, B => n1898, S => n2413, Z => n6251);
   U760 : MUX21L port map( A => n2482, B => n827, S => n2414, Z => n6250);
   U761 : MUX21L port map( A => n1897, B => n2482, S => n2415, Z => n6249);
   U762 : MUX21L port map( A => n826, B => n2482, S => n2416, Z => n6248);
   U763 : MUX21L port map( A => n1896, B => n2482, S => n2417, Z => n6247);
   U764 : MUX21L port map( A => n825, B => n2482, S => n2418, Z => n6246);
   U765 : MUX21L port map( A => n2482, B => n1903, S => n2419, Z => n6245);
   U766 : MUX21L port map( A => n2482, B => n832, S => n2420, Z => n6244);
   U767 : MUX21L port map( A => n2482, B => n1902, S => n2421, Z => n6243);
   U768 : MUX21L port map( A => n2482, B => n831, S => n2422, Z => n6242);
   U769 : MUX21L port map( A => n1901, B => n2482, S => n2423, Z => n6241);
   U770 : MUX21L port map( A => n830, B => n2482, S => n2424, Z => n6240);
   U771 : MUX21L port map( A => n1900, B => n2482, S => n2425, Z => n6239);
   U772 : MUX21L port map( A => n829, B => n2482, S => n2426, Z => n6238);
   U773 : MUX21L port map( A => n2482, B => n1907, S => n2427, Z => n6237);
   U774 : MUX21L port map( A => n2482, B => n836, S => n2428, Z => n6236);
   U775 : MUX21L port map( A => n2482, B => n1906, S => n2429, Z => n6235);
   U776 : MUX21L port map( A => n2482, B => n835, S => n2430, Z => n6234);
   U777 : MUX21L port map( A => n1905, B => n2482, S => n2431, Z => n6233);
   U778 : MUX21L port map( A => n834, B => n2482, S => n2432, Z => n6232);
   U779 : MUX21L port map( A => n1904, B => n2482, S => n2433, Z => n6231);
   U780 : MUX21L port map( A => n833, B => n2482, S => n2434, Z => n6230);
   U781 : MUX21L port map( A => n2482, B => n1911, S => n2435, Z => n6229);
   U782 : MUX21L port map( A => n2482, B => n840, S => n2436, Z => n6228);
   U783 : MUX21L port map( A => n2482, B => n1910, S => n2437, Z => n6227);
   U784 : MUX21L port map( A => n2482, B => n839, S => n2438, Z => n6226);
   U785 : MUX21L port map( A => n1909, B => n2482, S => n2439, Z => n6225);
   U786 : MUX21L port map( A => n838, B => n2482, S => n2440, Z => n6224);
   U787 : MUX21L port map( A => n1908, B => n2482, S => n2441, Z => n6223);
   U788 : MUX21L port map( A => n837, B => n2482, S => n2442, Z => n6222);
   U789 : MUX21L port map( A => n2482, B => n1883, S => n2443, Z => n6221);
   U790 : MUX21L port map( A => n2482, B => n812, S => n2444, Z => n6220);
   U791 : MUX21L port map( A => n2482, B => n1882, S => n2445, Z => n6219);
   U792 : MUX21L port map( A => n2482, B => n811, S => n2446, Z => n6218);
   U793 : MUX21L port map( A => n1881, B => n2482, S => n2447, Z => n6217);
   U794 : MUX21L port map( A => n810, B => n2482, S => n2448, Z => n6216);
   U795 : MUX21L port map( A => n1880, B => n2482, S => n2449, Z => n6215);
   U796 : MUX21L port map( A => n809, B => n2482, S => n2450, Z => n6214);
   U797 : MUX21L port map( A => n2482, B => n1887, S => n2451, Z => n6213);
   U798 : MUX21L port map( A => n2482, B => n816, S => n2452, Z => n6212);
   U799 : MUX21L port map( A => n2482, B => n1886, S => n2453, Z => n6211);
   U800 : MUX21L port map( A => n2482, B => n815, S => n2454, Z => n6210);
   U801 : MUX21L port map( A => n1885, B => n2482, S => n2455, Z => n6209);
   U802 : MUX21L port map( A => n814, B => n2482, S => n2456, Z => n6208);
   U803 : MUX21L port map( A => n1884, B => n2482, S => n2457, Z => n6207);
   U804 : MUX21L port map( A => n813, B => n2482, S => n2458, Z => n6206);
   U805 : MUX21L port map( A => n2482, B => n1891, S => n2459, Z => n6205);
   U806 : MUX21L port map( A => n2482, B => n820, S => n2460, Z => n6204);
   U807 : MUX21L port map( A => n2482, B => n1890, S => n2461, Z => n6203);
   U808 : MUX21L port map( A => n2482, B => n819, S => n2462, Z => n6202);
   U809 : MUX21L port map( A => n1889, B => n2482, S => n2463, Z => n6201);
   U810 : MUX21L port map( A => n818, B => n2482, S => n2464, Z => n6200);
   U811 : MUX21L port map( A => n1888, B => n2482, S => n2465, Z => n6199);
   U812 : MUX21L port map( A => n817, B => n2482, S => n2466, Z => n6198);
   U813 : MUX21L port map( A => n2482, B => n1895, S => n2467, Z => n6197);
   U814 : MUX21L port map( A => n2482, B => n824, S => n2468, Z => n6196);
   U815 : MUX21L port map( A => n2482, B => n1894, S => n2469, Z => n6195);
   U816 : MUX21L port map( A => n2482, B => n823, S => n2470, Z => n6194);
   U817 : MUX21L port map( A => n1893, B => n2482, S => n2471, Z => n6193);
   U818 : MUX21L port map( A => n822, B => n2482, S => n2472, Z => n6192);
   U819 : MUX21L port map( A => n1892, B => n2482, S => n2473, Z => n6191);
   U820 : MUX21L port map( A => n821, B => n2482, S => n2474, Z => n6190);
   U821 : AO2 port map( A => v_TEMP_VECTOR_25_port, B => n2475, C => 
                           v_KEY32_IN_25_port, D => n2476, Z => n2482);
   U822 : MUX21L port map( A => n2483, B => n2027, S => n2411, Z => n6189);
   U823 : MUX21L port map( A => n2483, B => n956, S => n2412, Z => n6188);
   U824 : MUX21L port map( A => n2483, B => n2026, S => n2413, Z => n6187);
   U825 : MUX21L port map( A => n2483, B => n955, S => n2414, Z => n6186);
   U826 : MUX21L port map( A => n2025, B => n2483, S => n2415, Z => n6185);
   U827 : MUX21L port map( A => n954, B => n2483, S => n2416, Z => n6184);
   U828 : MUX21L port map( A => n2024, B => n2483, S => n2417, Z => n6183);
   U829 : MUX21L port map( A => n953, B => n2483, S => n2418, Z => n6182);
   U830 : MUX21L port map( A => n2483, B => n2031, S => n2419, Z => n6181);
   U831 : MUX21L port map( A => n2483, B => n960, S => n2420, Z => n6180);
   U832 : MUX21L port map( A => n2483, B => n2030, S => n2421, Z => n6179);
   U833 : MUX21L port map( A => n2483, B => n959, S => n2422, Z => n6178);
   U834 : MUX21L port map( A => n2029, B => n2483, S => n2423, Z => n6177);
   U835 : MUX21L port map( A => n958, B => n2483, S => n2424, Z => n6176);
   U836 : MUX21L port map( A => n2028, B => n2483, S => n2425, Z => n6175);
   U837 : MUX21L port map( A => n957, B => n2483, S => n2426, Z => n6174);
   U838 : MUX21L port map( A => n2483, B => n2035, S => n2427, Z => n6173);
   U839 : MUX21L port map( A => n2483, B => n964, S => n2428, Z => n6172);
   U840 : MUX21L port map( A => n2483, B => n2034, S => n2429, Z => n6171);
   U841 : MUX21L port map( A => n2483, B => n963, S => n2430, Z => n6170);
   U842 : MUX21L port map( A => n2033, B => n2483, S => n2431, Z => n6169);
   U843 : MUX21L port map( A => n962, B => n2483, S => n2432, Z => n6168);
   U844 : MUX21L port map( A => n2032, B => n2483, S => n2433, Z => n6167);
   U845 : MUX21L port map( A => n961, B => n2483, S => n2434, Z => n6166);
   U846 : MUX21L port map( A => n2483, B => n2039, S => n2435, Z => n6165);
   U847 : MUX21L port map( A => n2483, B => n968, S => n2436, Z => n6164);
   U848 : MUX21L port map( A => n2483, B => n2038, S => n2437, Z => n6163);
   U849 : MUX21L port map( A => n2483, B => n967, S => n2438, Z => n6162);
   U850 : MUX21L port map( A => n2037, B => n2483, S => n2439, Z => n6161);
   U851 : MUX21L port map( A => n966, B => n2483, S => n2440, Z => n6160);
   U852 : MUX21L port map( A => n2036, B => n2483, S => n2441, Z => n6159);
   U853 : MUX21L port map( A => n965, B => n2483, S => n2442, Z => n6158);
   U854 : MUX21L port map( A => n2483, B => n2011, S => n2443, Z => n6157);
   U855 : MUX21L port map( A => n2483, B => n940, S => n2444, Z => n6156);
   U856 : MUX21L port map( A => n2483, B => n2010, S => n2445, Z => n6155);
   U857 : MUX21L port map( A => n2483, B => n939, S => n2446, Z => n6154);
   U858 : MUX21L port map( A => n2009, B => n2483, S => n2447, Z => n6153);
   U859 : MUX21L port map( A => n938, B => n2483, S => n2448, Z => n6152);
   U860 : MUX21L port map( A => n2008, B => n2483, S => n2449, Z => n6151);
   U861 : MUX21L port map( A => n937, B => n2483, S => n2450, Z => n6150);
   U862 : MUX21L port map( A => n2483, B => n2015, S => n2451, Z => n6149);
   U863 : MUX21L port map( A => n2483, B => n944, S => n2452, Z => n6148);
   U864 : MUX21L port map( A => n2483, B => n2014, S => n2453, Z => n6147);
   U865 : MUX21L port map( A => n2483, B => n943, S => n2454, Z => n6146);
   U866 : MUX21L port map( A => n2013, B => n2483, S => n2455, Z => n6145);
   U867 : MUX21L port map( A => n942, B => n2483, S => n2456, Z => n6144);
   U868 : MUX21L port map( A => n2012, B => n2483, S => n2457, Z => n6143);
   U869 : MUX21L port map( A => n941, B => n2483, S => n2458, Z => n6142);
   U870 : MUX21L port map( A => n2483, B => n2019, S => n2459, Z => n6141);
   U871 : MUX21L port map( A => n2483, B => n948, S => n2460, Z => n6140);
   U872 : MUX21L port map( A => n2483, B => n2018, S => n2461, Z => n6139);
   U873 : MUX21L port map( A => n2483, B => n947, S => n2462, Z => n6138);
   U874 : MUX21L port map( A => n2017, B => n2483, S => n2463, Z => n6137);
   U875 : MUX21L port map( A => n946, B => n2483, S => n2464, Z => n6136);
   U876 : MUX21L port map( A => n2016, B => n2483, S => n2465, Z => n6135);
   U877 : MUX21L port map( A => n945, B => n2483, S => n2466, Z => n6134);
   U878 : MUX21L port map( A => n2483, B => n2023, S => n2467, Z => n6133);
   U879 : MUX21L port map( A => n2483, B => n952, S => n2468, Z => n6132);
   U880 : MUX21L port map( A => n2483, B => n2022, S => n2469, Z => n6131);
   U881 : MUX21L port map( A => n2483, B => n951, S => n2470, Z => n6130);
   U882 : MUX21L port map( A => n2021, B => n2483, S => n2471, Z => n6129);
   U883 : MUX21L port map( A => n950, B => n2483, S => n2472, Z => n6128);
   U884 : MUX21L port map( A => n2020, B => n2483, S => n2473, Z => n6127);
   U885 : MUX21L port map( A => n949, B => n2483, S => n2474, Z => n6126);
   U886 : AO2 port map( A => v_TEMP_VECTOR_24_port, B => n2475, C => 
                           v_KEY32_IN_24_port, D => n2476, Z => n2483);
   U887 : MUX21L port map( A => n2484, B => n1163, S => n2411, Z => n6125);
   U888 : MUX21L port map( A => n2484, B => n92, S => n2412, Z => n6124);
   U889 : MUX21L port map( A => n2484, B => n1162, S => n2413, Z => n6123);
   U890 : MUX21L port map( A => n2484, B => n91, S => n2414, Z => n6122);
   U891 : MUX21L port map( A => n1161, B => n2484, S => n2415, Z => n6121);
   U892 : MUX21L port map( A => n90, B => n2484, S => n2416, Z => n6120);
   U893 : MUX21L port map( A => n1160, B => n2484, S => n2417, Z => n6119);
   U894 : MUX21L port map( A => n89, B => n2484, S => n2418, Z => n6118);
   U895 : MUX21L port map( A => n2484, B => n1167, S => n2419, Z => n6117);
   U896 : MUX21L port map( A => n2484, B => n96, S => n2420, Z => n6116);
   U897 : MUX21L port map( A => n2484, B => n1166, S => n2421, Z => n6115);
   U898 : MUX21L port map( A => n2484, B => n95, S => n2422, Z => n6114);
   U899 : MUX21L port map( A => n1165, B => n2484, S => n2423, Z => n6113);
   U900 : MUX21L port map( A => n94, B => n2484, S => n2424, Z => n6112);
   U901 : MUX21L port map( A => n1164, B => n2484, S => n2425, Z => n6111);
   U902 : MUX21L port map( A => n93, B => n2484, S => n2426, Z => n6110);
   U903 : MUX21L port map( A => n2484, B => n1171, S => n2427, Z => n6109);
   U904 : MUX21L port map( A => n2484, B => n100, S => n2428, Z => n6108);
   U905 : MUX21L port map( A => n2484, B => n1170, S => n2429, Z => n6107);
   U906 : MUX21L port map( A => n2484, B => n99, S => n2430, Z => n6106);
   U907 : MUX21L port map( A => n1169, B => n2484, S => n2431, Z => n6105);
   U908 : MUX21L port map( A => n98, B => n2484, S => n2432, Z => n6104);
   U909 : MUX21L port map( A => n1168, B => n2484, S => n2433, Z => n6103);
   U910 : MUX21L port map( A => n97, B => n2484, S => n2434, Z => n6102);
   U911 : MUX21L port map( A => n2484, B => n1175, S => n2435, Z => n6101);
   U912 : MUX21L port map( A => n2484, B => n104, S => n2436, Z => n6100);
   U913 : MUX21L port map( A => n2484, B => n1174, S => n2437, Z => n6099);
   U914 : MUX21L port map( A => n2484, B => n103, S => n2438, Z => n6098);
   U915 : MUX21L port map( A => n1173, B => n2484, S => n2439, Z => n6097);
   U916 : MUX21L port map( A => n102, B => n2484, S => n2440, Z => n6096);
   U917 : MUX21L port map( A => n1172, B => n2484, S => n2441, Z => n6095);
   U918 : MUX21L port map( A => n101, B => n2484, S => n2442, Z => n6094);
   U919 : MUX21L port map( A => n2484, B => n1147, S => n2443, Z => n6093);
   U920 : MUX21L port map( A => n2484, B => n76, S => n2444, Z => n6092);
   U921 : MUX21L port map( A => n2484, B => n1146, S => n2445, Z => n6091);
   U922 : MUX21L port map( A => n2484, B => n75, S => n2446, Z => n6090);
   U923 : MUX21L port map( A => n1145, B => n2484, S => n2447, Z => n6089);
   U924 : MUX21L port map( A => n74, B => n2484, S => n2448, Z => n6088);
   U925 : MUX21L port map( A => n1144, B => n2484, S => n2449, Z => n6087);
   U926 : MUX21L port map( A => n73, B => n2484, S => n2450, Z => n6086);
   U927 : MUX21L port map( A => n2484, B => n1151, S => n2451, Z => n6085);
   U928 : MUX21L port map( A => n2484, B => n80, S => n2452, Z => n6084);
   U929 : MUX21L port map( A => n2484, B => n1150, S => n2453, Z => n6083);
   U930 : MUX21L port map( A => n2484, B => n79, S => n2454, Z => n6082);
   U931 : MUX21L port map( A => n1149, B => n2484, S => n2455, Z => n6081);
   U932 : MUX21L port map( A => n78, B => n2484, S => n2456, Z => n6080);
   U933 : MUX21L port map( A => n1148, B => n2484, S => n2457, Z => n6079);
   U934 : MUX21L port map( A => n77, B => n2484, S => n2458, Z => n6078);
   U935 : MUX21L port map( A => n2484, B => n1155, S => n2459, Z => n6077);
   U936 : MUX21L port map( A => n2484, B => n84, S => n2460, Z => n6076);
   U937 : MUX21L port map( A => n2484, B => n1154, S => n2461, Z => n6075);
   U938 : MUX21L port map( A => n2484, B => n83, S => n2462, Z => n6074);
   U939 : MUX21L port map( A => n1153, B => n2484, S => n2463, Z => n6073);
   U940 : MUX21L port map( A => n82, B => n2484, S => n2464, Z => n6072);
   U941 : MUX21L port map( A => n1152, B => n2484, S => n2465, Z => n6071);
   U942 : MUX21L port map( A => n81, B => n2484, S => n2466, Z => n6070);
   U943 : MUX21L port map( A => n2484, B => n1159, S => n2467, Z => n6069);
   U944 : MUX21L port map( A => n2484, B => n88, S => n2468, Z => n6068);
   U945 : MUX21L port map( A => n2484, B => n1158, S => n2469, Z => n6067);
   U946 : MUX21L port map( A => n2484, B => n87, S => n2470, Z => n6066);
   U947 : MUX21L port map( A => n1157, B => n2484, S => n2471, Z => n6065);
   U948 : MUX21L port map( A => n86, B => n2484, S => n2472, Z => n6064);
   U949 : MUX21L port map( A => n1156, B => n2484, S => n2473, Z => n6063);
   U950 : MUX21L port map( A => n85, B => n2484, S => n2474, Z => n6062);
   U951 : AO2 port map( A => v_TEMP_VECTOR_23_port, B => n2475, C => 
                           v_KEY32_IN_23_port, D => n2476, Z => n2484);
   U952 : MUX21L port map( A => n2485, B => n1291, S => n2411, Z => n6061);
   U953 : MUX21L port map( A => n2485, B => n220, S => n2412, Z => n6060);
   U954 : MUX21L port map( A => n2485, B => n1290, S => n2413, Z => n6059);
   U955 : MUX21L port map( A => n2485, B => n219, S => n2414, Z => n6058);
   U956 : MUX21L port map( A => n1289, B => n2485, S => n2415, Z => n6057);
   U957 : MUX21L port map( A => n218, B => n2485, S => n2416, Z => n6056);
   U958 : MUX21L port map( A => n1288, B => n2485, S => n2417, Z => n6055);
   U959 : MUX21L port map( A => n217, B => n2485, S => n2418, Z => n6054);
   U960 : MUX21L port map( A => n2485, B => n1295, S => n2419, Z => n6053);
   U961 : MUX21L port map( A => n2485, B => n224, S => n2420, Z => n6052);
   U962 : MUX21L port map( A => n2485, B => n1294, S => n2421, Z => n6051);
   U963 : MUX21L port map( A => n2485, B => n223, S => n2422, Z => n6050);
   U964 : MUX21L port map( A => n1293, B => n2485, S => n2423, Z => n6049);
   U965 : MUX21L port map( A => n222, B => n2485, S => n2424, Z => n6048);
   U966 : MUX21L port map( A => n1292, B => n2485, S => n2425, Z => n6047);
   U967 : MUX21L port map( A => n221, B => n2485, S => n2426, Z => n6046);
   U968 : MUX21L port map( A => n2485, B => n1299, S => n2427, Z => n6045);
   U969 : MUX21L port map( A => n2485, B => n228, S => n2428, Z => n6044);
   U970 : MUX21L port map( A => n2485, B => n1298, S => n2429, Z => n6043);
   U971 : MUX21L port map( A => n2485, B => n227, S => n2430, Z => n6042);
   U972 : MUX21L port map( A => n1297, B => n2485, S => n2431, Z => n6041);
   U973 : MUX21L port map( A => n226, B => n2485, S => n2432, Z => n6040);
   U974 : MUX21L port map( A => n1296, B => n2485, S => n2433, Z => n6039);
   U975 : MUX21L port map( A => n225, B => n2485, S => n2434, Z => n6038);
   U976 : MUX21L port map( A => n2485, B => n1303, S => n2435, Z => n6037);
   U977 : MUX21L port map( A => n2485, B => n232, S => n2436, Z => n6036);
   U978 : MUX21L port map( A => n2485, B => n1302, S => n2437, Z => n6035);
   U979 : MUX21L port map( A => n2485, B => n231, S => n2438, Z => n6034);
   U980 : MUX21L port map( A => n1301, B => n2485, S => n2439, Z => n6033);
   U981 : MUX21L port map( A => n230, B => n2485, S => n2440, Z => n6032);
   U982 : MUX21L port map( A => n1300, B => n2485, S => n2441, Z => n6031);
   U983 : MUX21L port map( A => n229, B => n2485, S => n2442, Z => n6030);
   U984 : MUX21L port map( A => n2485, B => n1275, S => n2443, Z => n6029);
   U985 : MUX21L port map( A => n2485, B => n204, S => n2444, Z => n6028);
   U986 : MUX21L port map( A => n2485, B => n1274, S => n2445, Z => n6027);
   U987 : MUX21L port map( A => n2485, B => n203, S => n2446, Z => n6026);
   U988 : MUX21L port map( A => n1273, B => n2485, S => n2447, Z => n6025);
   U989 : MUX21L port map( A => n202, B => n2485, S => n2448, Z => n6024);
   U990 : MUX21L port map( A => n1272, B => n2485, S => n2449, Z => n6023);
   U991 : MUX21L port map( A => n201, B => n2485, S => n2450, Z => n6022);
   U992 : MUX21L port map( A => n2485, B => n1279, S => n2451, Z => n6021);
   U993 : MUX21L port map( A => n2485, B => n208, S => n2452, Z => n6020);
   U994 : MUX21L port map( A => n2485, B => n1278, S => n2453, Z => n6019);
   U995 : MUX21L port map( A => n2485, B => n207, S => n2454, Z => n6018);
   U996 : MUX21L port map( A => n1277, B => n2485, S => n2455, Z => n6017);
   U997 : MUX21L port map( A => n206, B => n2485, S => n2456, Z => n6016);
   U998 : MUX21L port map( A => n1276, B => n2485, S => n2457, Z => n6015);
   U999 : MUX21L port map( A => n205, B => n2485, S => n2458, Z => n6014);
   U1000 : MUX21L port map( A => n2485, B => n1283, S => n2459, Z => n6013);
   U1001 : MUX21L port map( A => n2485, B => n212, S => n2460, Z => n6012);
   U1002 : MUX21L port map( A => n2485, B => n1282, S => n2461, Z => n6011);
   U1003 : MUX21L port map( A => n2485, B => n211, S => n2462, Z => n6010);
   U1004 : MUX21L port map( A => n1281, B => n2485, S => n2463, Z => n6009);
   U1005 : MUX21L port map( A => n210, B => n2485, S => n2464, Z => n6008);
   U1006 : MUX21L port map( A => n1280, B => n2485, S => n2465, Z => n6007);
   U1007 : MUX21L port map( A => n209, B => n2485, S => n2466, Z => n6006);
   U1008 : MUX21L port map( A => n2485, B => n1287, S => n2467, Z => n6005);
   U1009 : MUX21L port map( A => n2485, B => n216, S => n2468, Z => n6004);
   U1010 : MUX21L port map( A => n2485, B => n1286, S => n2469, Z => n6003);
   U1011 : MUX21L port map( A => n2485, B => n215, S => n2470, Z => n6002);
   U1012 : MUX21L port map( A => n1285, B => n2485, S => n2471, Z => n6001);
   U1013 : MUX21L port map( A => n214, B => n2485, S => n2472, Z => n6000);
   U1014 : MUX21L port map( A => n1284, B => n2485, S => n2473, Z => n5999);
   U1015 : MUX21L port map( A => n213, B => n2485, S => n2474, Z => n5998);
   U1016 : AO2 port map( A => v_TEMP_VECTOR_22_port, B => n2475, C => 
                           v_KEY32_IN_22_port, D => n2476, Z => n2485);
   U1017 : MUX21L port map( A => n2486, B => n1419, S => n2411, Z => n5997);
   U1018 : MUX21L port map( A => n2486, B => n348, S => n2412, Z => n5996);
   U1019 : MUX21L port map( A => n2486, B => n1418, S => n2413, Z => n5995);
   U1020 : MUX21L port map( A => n2486, B => n347, S => n2414, Z => n5994);
   U1021 : MUX21L port map( A => n1417, B => n2486, S => n2415, Z => n5993);
   U1022 : MUX21L port map( A => n346, B => n2486, S => n2416, Z => n5992);
   U1023 : MUX21L port map( A => n1416, B => n2486, S => n2417, Z => n5991);
   U1024 : MUX21L port map( A => n345, B => n2486, S => n2418, Z => n5990);
   U1025 : MUX21L port map( A => n2486, B => n1423, S => n2419, Z => n5989);
   U1026 : MUX21L port map( A => n2486, B => n352, S => n2420, Z => n5988);
   U1027 : MUX21L port map( A => n2486, B => n1422, S => n2421, Z => n5987);
   U1028 : MUX21L port map( A => n2486, B => n351, S => n2422, Z => n5986);
   U1029 : MUX21L port map( A => n1421, B => n2486, S => n2423, Z => n5985);
   U1030 : MUX21L port map( A => n350, B => n2486, S => n2424, Z => n5984);
   U1031 : MUX21L port map( A => n1420, B => n2486, S => n2425, Z => n5983);
   U1032 : MUX21L port map( A => n349, B => n2486, S => n2426, Z => n5982);
   U1033 : MUX21L port map( A => n2486, B => n1427, S => n2427, Z => n5981);
   U1034 : MUX21L port map( A => n2486, B => n356, S => n2428, Z => n5980);
   U1035 : MUX21L port map( A => n2486, B => n1426, S => n2429, Z => n5979);
   U1036 : MUX21L port map( A => n2486, B => n355, S => n2430, Z => n5978);
   U1037 : MUX21L port map( A => n1425, B => n2486, S => n2431, Z => n5977);
   U1038 : MUX21L port map( A => n354, B => n2486, S => n2432, Z => n5976);
   U1039 : MUX21L port map( A => n1424, B => n2486, S => n2433, Z => n5975);
   U1040 : MUX21L port map( A => n353, B => n2486, S => n2434, Z => n5974);
   U1041 : MUX21L port map( A => n2486, B => n1431, S => n2435, Z => n5973);
   U1042 : MUX21L port map( A => n2486, B => n360, S => n2436, Z => n5972);
   U1043 : MUX21L port map( A => n2486, B => n1430, S => n2437, Z => n5971);
   U1044 : MUX21L port map( A => n2486, B => n359, S => n2438, Z => n5970);
   U1045 : MUX21L port map( A => n1429, B => n2486, S => n2439, Z => n5969);
   U1046 : MUX21L port map( A => n358, B => n2486, S => n2440, Z => n5968);
   U1047 : MUX21L port map( A => n1428, B => n2486, S => n2441, Z => n5967);
   U1048 : MUX21L port map( A => n357, B => n2486, S => n2442, Z => n5966);
   U1049 : MUX21L port map( A => n2486, B => n1403, S => n2443, Z => n5965);
   U1050 : MUX21L port map( A => n2486, B => n332, S => n2444, Z => n5964);
   U1051 : MUX21L port map( A => n2486, B => n1402, S => n2445, Z => n5963);
   U1052 : MUX21L port map( A => n2486, B => n331, S => n2446, Z => n5962);
   U1053 : MUX21L port map( A => n1401, B => n2486, S => n2447, Z => n5961);
   U1054 : MUX21L port map( A => n330, B => n2486, S => n2448, Z => n5960);
   U1055 : MUX21L port map( A => n1400, B => n2486, S => n2449, Z => n5959);
   U1056 : MUX21L port map( A => n329, B => n2486, S => n2450, Z => n5958);
   U1057 : MUX21L port map( A => n2486, B => n1407, S => n2451, Z => n5957);
   U1058 : MUX21L port map( A => n2486, B => n336, S => n2452, Z => n5956);
   U1059 : MUX21L port map( A => n2486, B => n1406, S => n2453, Z => n5955);
   U1060 : MUX21L port map( A => n2486, B => n335, S => n2454, Z => n5954);
   U1061 : MUX21L port map( A => n1405, B => n2486, S => n2455, Z => n5953);
   U1062 : MUX21L port map( A => n334, B => n2486, S => n2456, Z => n5952);
   U1063 : MUX21L port map( A => n1404, B => n2486, S => n2457, Z => n5951);
   U1064 : MUX21L port map( A => n333, B => n2486, S => n2458, Z => n5950);
   U1065 : MUX21L port map( A => n2486, B => n1411, S => n2459, Z => n5949);
   U1066 : MUX21L port map( A => n2486, B => n340, S => n2460, Z => n5948);
   U1067 : MUX21L port map( A => n2486, B => n1410, S => n2461, Z => n5947);
   U1068 : MUX21L port map( A => n2486, B => n339, S => n2462, Z => n5946);
   U1069 : MUX21L port map( A => n1409, B => n2486, S => n2463, Z => n5945);
   U1070 : MUX21L port map( A => n338, B => n2486, S => n2464, Z => n5944);
   U1071 : MUX21L port map( A => n1408, B => n2486, S => n2465, Z => n5943);
   U1072 : MUX21L port map( A => n337, B => n2486, S => n2466, Z => n5942);
   U1073 : MUX21L port map( A => n2486, B => n1415, S => n2467, Z => n5941);
   U1074 : MUX21L port map( A => n2486, B => n344, S => n2468, Z => n5940);
   U1075 : MUX21L port map( A => n2486, B => n1414, S => n2469, Z => n5939);
   U1076 : MUX21L port map( A => n2486, B => n343, S => n2470, Z => n5938);
   U1077 : MUX21L port map( A => n1413, B => n2486, S => n2471, Z => n5937);
   U1078 : MUX21L port map( A => n342, B => n2486, S => n2472, Z => n5936);
   U1079 : MUX21L port map( A => n1412, B => n2486, S => n2473, Z => n5935);
   U1080 : MUX21L port map( A => n341, B => n2486, S => n2474, Z => n5934);
   U1081 : AO2 port map( A => v_TEMP_VECTOR_21_port, B => n2475, C => 
                           v_KEY32_IN_21_port, D => n2476, Z => n2486);
   U1082 : MUX21L port map( A => n2487, B => n1547, S => n2411, Z => n5933);
   U1083 : MUX21L port map( A => n2487, B => n476, S => n2412, Z => n5932);
   U1084 : MUX21L port map( A => n2487, B => n1546, S => n2413, Z => n5931);
   U1085 : MUX21L port map( A => n2487, B => n475, S => n2414, Z => n5930);
   U1086 : MUX21L port map( A => n1545, B => n2487, S => n2415, Z => n5929);
   U1087 : MUX21L port map( A => n474, B => n2487, S => n2416, Z => n5928);
   U1088 : MUX21L port map( A => n1544, B => n2487, S => n2417, Z => n5927);
   U1089 : MUX21L port map( A => n473, B => n2487, S => n2418, Z => n5926);
   U1090 : MUX21L port map( A => n2487, B => n1551, S => n2419, Z => n5925);
   U1091 : MUX21L port map( A => n2487, B => n480, S => n2420, Z => n5924);
   U1092 : MUX21L port map( A => n2487, B => n1550, S => n2421, Z => n5923);
   U1093 : MUX21L port map( A => n2487, B => n479, S => n2422, Z => n5922);
   U1094 : MUX21L port map( A => n1549, B => n2487, S => n2423, Z => n5921);
   U1095 : MUX21L port map( A => n478, B => n2487, S => n2424, Z => n5920);
   U1096 : MUX21L port map( A => n1548, B => n2487, S => n2425, Z => n5919);
   U1097 : MUX21L port map( A => n477, B => n2487, S => n2426, Z => n5918);
   U1098 : MUX21L port map( A => n2487, B => n1555, S => n2427, Z => n5917);
   U1099 : MUX21L port map( A => n2487, B => n484, S => n2428, Z => n5916);
   U1100 : MUX21L port map( A => n2487, B => n1554, S => n2429, Z => n5915);
   U1101 : MUX21L port map( A => n2487, B => n483, S => n2430, Z => n5914);
   U1102 : MUX21L port map( A => n1553, B => n2487, S => n2431, Z => n5913);
   U1103 : MUX21L port map( A => n482, B => n2487, S => n2432, Z => n5912);
   U1104 : MUX21L port map( A => n1552, B => n2487, S => n2433, Z => n5911);
   U1105 : MUX21L port map( A => n481, B => n2487, S => n2434, Z => n5910);
   U1106 : MUX21L port map( A => n2487, B => n1559, S => n2435, Z => n5909);
   U1107 : MUX21L port map( A => n2487, B => n488, S => n2436, Z => n5908);
   U1108 : MUX21L port map( A => n2487, B => n1558, S => n2437, Z => n5907);
   U1109 : MUX21L port map( A => n2487, B => n487, S => n2438, Z => n5906);
   U1110 : MUX21L port map( A => n1557, B => n2487, S => n2439, Z => n5905);
   U1111 : MUX21L port map( A => n486, B => n2487, S => n2440, Z => n5904);
   U1112 : MUX21L port map( A => n1556, B => n2487, S => n2441, Z => n5903);
   U1113 : MUX21L port map( A => n485, B => n2487, S => n2442, Z => n5902);
   U1114 : MUX21L port map( A => n2487, B => n1531, S => n2443, Z => n5901);
   U1115 : MUX21L port map( A => n2487, B => n460, S => n2444, Z => n5900);
   U1116 : MUX21L port map( A => n2487, B => n1530, S => n2445, Z => n5899);
   U1117 : MUX21L port map( A => n2487, B => n459, S => n2446, Z => n5898);
   U1118 : MUX21L port map( A => n1529, B => n2487, S => n2447, Z => n5897);
   U1119 : MUX21L port map( A => n458, B => n2487, S => n2448, Z => n5896);
   U1120 : MUX21L port map( A => n1528, B => n2487, S => n2449, Z => n5895);
   U1121 : MUX21L port map( A => n457, B => n2487, S => n2450, Z => n5894);
   U1122 : MUX21L port map( A => n2487, B => n1535, S => n2451, Z => n5893);
   U1123 : MUX21L port map( A => n2487, B => n464, S => n2452, Z => n5892);
   U1124 : MUX21L port map( A => n2487, B => n1534, S => n2453, Z => n5891);
   U1125 : MUX21L port map( A => n2487, B => n463, S => n2454, Z => n5890);
   U1126 : MUX21L port map( A => n1533, B => n2487, S => n2455, Z => n5889);
   U1127 : MUX21L port map( A => n462, B => n2487, S => n2456, Z => n5888);
   U1128 : MUX21L port map( A => n1532, B => n2487, S => n2457, Z => n5887);
   U1129 : MUX21L port map( A => n461, B => n2487, S => n2458, Z => n5886);
   U1130 : MUX21L port map( A => n2487, B => n1539, S => n2459, Z => n5885);
   U1131 : MUX21L port map( A => n2487, B => n468, S => n2460, Z => n5884);
   U1132 : MUX21L port map( A => n2487, B => n1538, S => n2461, Z => n5883);
   U1133 : MUX21L port map( A => n2487, B => n467, S => n2462, Z => n5882);
   U1134 : MUX21L port map( A => n1537, B => n2487, S => n2463, Z => n5881);
   U1135 : MUX21L port map( A => n466, B => n2487, S => n2464, Z => n5880);
   U1136 : MUX21L port map( A => n1536, B => n2487, S => n2465, Z => n5879);
   U1137 : MUX21L port map( A => n465, B => n2487, S => n2466, Z => n5878);
   U1138 : MUX21L port map( A => n2487, B => n1543, S => n2467, Z => n5877);
   U1139 : MUX21L port map( A => n2487, B => n472, S => n2468, Z => n5876);
   U1140 : MUX21L port map( A => n2487, B => n1542, S => n2469, Z => n5875);
   U1141 : MUX21L port map( A => n2487, B => n471, S => n2470, Z => n5874);
   U1142 : MUX21L port map( A => n1541, B => n2487, S => n2471, Z => n5873);
   U1143 : MUX21L port map( A => n470, B => n2487, S => n2472, Z => n5872);
   U1144 : MUX21L port map( A => n1540, B => n2487, S => n2473, Z => n5871);
   U1145 : MUX21L port map( A => n469, B => n2487, S => n2474, Z => n5870);
   U1146 : AO2 port map( A => v_TEMP_VECTOR_20_port, B => n2475, C => 
                           v_KEY32_IN_20_port, D => n2476, Z => n2487);
   U1147 : MUX21L port map( A => n2488, B => n1675, S => n2411, Z => n5869);
   U1148 : MUX21L port map( A => n2488, B => n604, S => n2412, Z => n5868);
   U1149 : MUX21L port map( A => n2488, B => n1674, S => n2413, Z => n5867);
   U1150 : MUX21L port map( A => n2488, B => n603, S => n2414, Z => n5866);
   U1151 : MUX21L port map( A => n1673, B => n2488, S => n2415, Z => n5865);
   U1152 : MUX21L port map( A => n602, B => n2488, S => n2416, Z => n5864);
   U1153 : MUX21L port map( A => n1672, B => n2488, S => n2417, Z => n5863);
   U1154 : MUX21L port map( A => n601, B => n2488, S => n2418, Z => n5862);
   U1155 : MUX21L port map( A => n2488, B => n1679, S => n2419, Z => n5861);
   U1156 : MUX21L port map( A => n2488, B => n608, S => n2420, Z => n5860);
   U1157 : MUX21L port map( A => n2488, B => n1678, S => n2421, Z => n5859);
   U1158 : MUX21L port map( A => n2488, B => n607, S => n2422, Z => n5858);
   U1159 : MUX21L port map( A => n1677, B => n2488, S => n2423, Z => n5857);
   U1160 : MUX21L port map( A => n606, B => n2488, S => n2424, Z => n5856);
   U1161 : MUX21L port map( A => n1676, B => n2488, S => n2425, Z => n5855);
   U1162 : MUX21L port map( A => n605, B => n2488, S => n2426, Z => n5854);
   U1163 : MUX21L port map( A => n2488, B => n1683, S => n2427, Z => n5853);
   U1164 : MUX21L port map( A => n2488, B => n612, S => n2428, Z => n5852);
   U1165 : MUX21L port map( A => n2488, B => n1682, S => n2429, Z => n5851);
   U1166 : MUX21L port map( A => n2488, B => n611, S => n2430, Z => n5850);
   U1167 : MUX21L port map( A => n1681, B => n2488, S => n2431, Z => n5849);
   U1168 : MUX21L port map( A => n610, B => n2488, S => n2432, Z => n5848);
   U1169 : MUX21L port map( A => n1680, B => n2488, S => n2433, Z => n5847);
   U1170 : MUX21L port map( A => n609, B => n2488, S => n2434, Z => n5846);
   U1171 : MUX21L port map( A => n2488, B => n1687, S => n2435, Z => n5845);
   U1172 : MUX21L port map( A => n2488, B => n616, S => n2436, Z => n5844);
   U1173 : MUX21L port map( A => n2488, B => n1686, S => n2437, Z => n5843);
   U1174 : MUX21L port map( A => n2488, B => n615, S => n2438, Z => n5842);
   U1175 : MUX21L port map( A => n1685, B => n2488, S => n2439, Z => n5841);
   U1176 : MUX21L port map( A => n614, B => n2488, S => n2440, Z => n5840);
   U1177 : MUX21L port map( A => n1684, B => n2488, S => n2441, Z => n5839);
   U1178 : MUX21L port map( A => n613, B => n2488, S => n2442, Z => n5838);
   U1179 : MUX21L port map( A => n2488, B => n1659, S => n2443, Z => n5837);
   U1180 : MUX21L port map( A => n2488, B => n588, S => n2444, Z => n5836);
   U1181 : MUX21L port map( A => n2488, B => n1658, S => n2445, Z => n5835);
   U1182 : MUX21L port map( A => n2488, B => n587, S => n2446, Z => n5834);
   U1183 : MUX21L port map( A => n1657, B => n2488, S => n2447, Z => n5833);
   U1184 : MUX21L port map( A => n586, B => n2488, S => n2448, Z => n5832);
   U1185 : MUX21L port map( A => n1656, B => n2488, S => n2449, Z => n5831);
   U1186 : MUX21L port map( A => n585, B => n2488, S => n2450, Z => n5830);
   U1187 : MUX21L port map( A => n2488, B => n1663, S => n2451, Z => n5829);
   U1188 : MUX21L port map( A => n2488, B => n592, S => n2452, Z => n5828);
   U1189 : MUX21L port map( A => n2488, B => n1662, S => n2453, Z => n5827);
   U1190 : MUX21L port map( A => n2488, B => n591, S => n2454, Z => n5826);
   U1191 : MUX21L port map( A => n1661, B => n2488, S => n2455, Z => n5825);
   U1192 : MUX21L port map( A => n590, B => n2488, S => n2456, Z => n5824);
   U1193 : MUX21L port map( A => n1660, B => n2488, S => n2457, Z => n5823);
   U1194 : MUX21L port map( A => n589, B => n2488, S => n2458, Z => n5822);
   U1195 : MUX21L port map( A => n2488, B => n1667, S => n2459, Z => n5821);
   U1196 : MUX21L port map( A => n2488, B => n596, S => n2460, Z => n5820);
   U1197 : MUX21L port map( A => n2488, B => n1666, S => n2461, Z => n5819);
   U1198 : MUX21L port map( A => n2488, B => n595, S => n2462, Z => n5818);
   U1199 : MUX21L port map( A => n1665, B => n2488, S => n2463, Z => n5817);
   U1200 : MUX21L port map( A => n594, B => n2488, S => n2464, Z => n5816);
   U1201 : MUX21L port map( A => n1664, B => n2488, S => n2465, Z => n5815);
   U1202 : MUX21L port map( A => n593, B => n2488, S => n2466, Z => n5814);
   U1203 : MUX21L port map( A => n2488, B => n1671, S => n2467, Z => n5813);
   U1204 : MUX21L port map( A => n2488, B => n600, S => n2468, Z => n5812);
   U1205 : MUX21L port map( A => n2488, B => n1670, S => n2469, Z => n5811);
   U1206 : MUX21L port map( A => n2488, B => n599, S => n2470, Z => n5810);
   U1207 : MUX21L port map( A => n1669, B => n2488, S => n2471, Z => n5809);
   U1208 : MUX21L port map( A => n598, B => n2488, S => n2472, Z => n5808);
   U1209 : MUX21L port map( A => n1668, B => n2488, S => n2473, Z => n5807);
   U1210 : MUX21L port map( A => n597, B => n2488, S => n2474, Z => n5806);
   U1211 : AO2 port map( A => v_TEMP_VECTOR_19_port, B => n2475, C => 
                           v_KEY32_IN_19_port, D => n2476, Z => n2488);
   U1212 : MUX21L port map( A => n2490, B => n1803, S => n2411, Z => n5805);
   U1213 : MUX21L port map( A => n2490, B => n732, S => n2412, Z => n5804);
   U1214 : MUX21L port map( A => n2490, B => n1802, S => n2413, Z => n5803);
   U1215 : MUX21L port map( A => n2490, B => n731, S => n2414, Z => n5802);
   U1216 : MUX21L port map( A => n1801, B => n2490, S => n2415, Z => n5801);
   U1217 : MUX21L port map( A => n730, B => n2490, S => n2416, Z => n5800);
   U1218 : MUX21L port map( A => n1800, B => n2490, S => n2417, Z => n5799);
   U1219 : MUX21L port map( A => n729, B => n2490, S => n2418, Z => n5798);
   U1220 : MUX21L port map( A => n2490, B => n1807, S => n2419, Z => n5797);
   U1221 : MUX21L port map( A => n2490, B => n736, S => n2420, Z => n5796);
   U1222 : MUX21L port map( A => n2490, B => n1806, S => n2421, Z => n5795);
   U1223 : MUX21L port map( A => n2490, B => n735, S => n2422, Z => n5794);
   U1224 : MUX21L port map( A => n1805, B => n2490, S => n2423, Z => n5793);
   U1225 : MUX21L port map( A => n734, B => n2490, S => n2424, Z => n5792);
   U1226 : MUX21L port map( A => n1804, B => n2490, S => n2425, Z => n5791);
   U1227 : MUX21L port map( A => n733, B => n2490, S => n2426, Z => n5790);
   U1228 : MUX21L port map( A => n2490, B => n1811, S => n2427, Z => n5789);
   U1229 : MUX21L port map( A => n2490, B => n740, S => n2428, Z => n5788);
   U1230 : MUX21L port map( A => n2490, B => n1810, S => n2429, Z => n5787);
   U1231 : MUX21L port map( A => n2490, B => n739, S => n2430, Z => n5786);
   U1232 : MUX21L port map( A => n1809, B => n2490, S => n2431, Z => n5785);
   U1233 : MUX21L port map( A => n738, B => n2490, S => n2432, Z => n5784);
   U1234 : MUX21L port map( A => n1808, B => n2490, S => n2433, Z => n5783);
   U1235 : MUX21L port map( A => n737, B => n2490, S => n2434, Z => n5782);
   U1236 : MUX21L port map( A => n2490, B => n1815, S => n2435, Z => n5781);
   U1237 : MUX21L port map( A => n2490, B => n744, S => n2436, Z => n5780);
   U1238 : MUX21L port map( A => n2490, B => n1814, S => n2437, Z => n5779);
   U1239 : MUX21L port map( A => n2490, B => n743, S => n2438, Z => n5778);
   U1240 : MUX21L port map( A => n1813, B => n2490, S => n2439, Z => n5777);
   U1241 : MUX21L port map( A => n742, B => n2490, S => n2440, Z => n5776);
   U1242 : MUX21L port map( A => n1812, B => n2490, S => n2441, Z => n5775);
   U1243 : MUX21L port map( A => n741, B => n2490, S => n2442, Z => n5774);
   U1244 : MUX21L port map( A => n2490, B => n1787, S => n2443, Z => n5773);
   U1245 : MUX21L port map( A => n2490, B => n716, S => n2444, Z => n5772);
   U1246 : MUX21L port map( A => n2490, B => n1786, S => n2445, Z => n5771);
   U1247 : MUX21L port map( A => n2490, B => n715, S => n2446, Z => n5770);
   U1248 : MUX21L port map( A => n1785, B => n2490, S => n2447, Z => n5769);
   U1249 : MUX21L port map( A => n714, B => n2490, S => n2448, Z => n5768);
   U1250 : MUX21L port map( A => n1784, B => n2490, S => n2449, Z => n5767);
   U1251 : MUX21L port map( A => n713, B => n2490, S => n2450, Z => n5766);
   U1252 : MUX21L port map( A => n2490, B => n1791, S => n2451, Z => n5765);
   U1253 : MUX21L port map( A => n2490, B => n720, S => n2452, Z => n5764);
   U1254 : MUX21L port map( A => n2490, B => n1790, S => n2453, Z => n5763);
   U1255 : MUX21L port map( A => n2490, B => n719, S => n2454, Z => n5762);
   U1256 : MUX21L port map( A => n1789, B => n2490, S => n2455, Z => n5761);
   U1257 : MUX21L port map( A => n718, B => n2490, S => n2456, Z => n5760);
   U1258 : MUX21L port map( A => n1788, B => n2490, S => n2457, Z => n5759);
   U1259 : MUX21L port map( A => n717, B => n2490, S => n2458, Z => n5758);
   U1260 : MUX21L port map( A => n2490, B => n1795, S => n2459, Z => n5757);
   U1261 : MUX21L port map( A => n2490, B => n724, S => n2460, Z => n5756);
   U1262 : MUX21L port map( A => n2490, B => n1794, S => n2461, Z => n5755);
   U1263 : MUX21L port map( A => n2490, B => n723, S => n2462, Z => n5754);
   U1264 : MUX21L port map( A => n1793, B => n2490, S => n2463, Z => n5753);
   U1265 : MUX21L port map( A => n722, B => n2490, S => n2464, Z => n5752);
   U1266 : MUX21L port map( A => n1792, B => n2490, S => n2465, Z => n5751);
   U1267 : MUX21L port map( A => n721, B => n2490, S => n2466, Z => n5750);
   U1268 : MUX21L port map( A => n2490, B => n1799, S => n2467, Z => n5749);
   U1269 : MUX21L port map( A => n2490, B => n728, S => n2468, Z => n5748);
   U1270 : MUX21L port map( A => n2490, B => n1798, S => n2469, Z => n5747);
   U1271 : MUX21L port map( A => n2490, B => n727, S => n2470, Z => n5746);
   U1272 : MUX21L port map( A => n1797, B => n2490, S => n2471, Z => n5745);
   U1273 : MUX21L port map( A => n726, B => n2490, S => n2472, Z => n5744);
   U1274 : MUX21L port map( A => n1796, B => n2490, S => n2473, Z => n5743);
   U1275 : MUX21L port map( A => n725, B => n2490, S => n2474, Z => n5742);
   U1276 : AO2 port map( A => v_TEMP_VECTOR_18_port, B => n2475, C => 
                           v_KEY32_IN_18_port, D => n2476, Z => n2490);
   U1277 : MUX21L port map( A => n2491, B => n1931, S => n2411, Z => n5741);
   U1278 : MUX21L port map( A => n2491, B => n860, S => n2412, Z => n5740);
   U1279 : MUX21L port map( A => n2491, B => n1930, S => n2413, Z => n5739);
   U1280 : MUX21L port map( A => n2491, B => n859, S => n2414, Z => n5738);
   U1281 : MUX21L port map( A => n1929, B => n2491, S => n2415, Z => n5737);
   U1282 : MUX21L port map( A => n858, B => n2491, S => n2416, Z => n5736);
   U1283 : MUX21L port map( A => n1928, B => n2491, S => n2417, Z => n5735);
   U1284 : MUX21L port map( A => n857, B => n2491, S => n2418, Z => n5734);
   U1285 : MUX21L port map( A => n2491, B => n1935, S => n2419, Z => n5733);
   U1286 : MUX21L port map( A => n2491, B => n864, S => n2420, Z => n5732);
   U1287 : MUX21L port map( A => n2491, B => n1934, S => n2421, Z => n5731);
   U1288 : MUX21L port map( A => n2491, B => n863, S => n2422, Z => n5730);
   U1289 : MUX21L port map( A => n1933, B => n2491, S => n2423, Z => n5729);
   U1290 : MUX21L port map( A => n862, B => n2491, S => n2424, Z => n5728);
   U1291 : MUX21L port map( A => n1932, B => n2491, S => n2425, Z => n5727);
   U1292 : MUX21L port map( A => n861, B => n2491, S => n2426, Z => n5726);
   U1293 : MUX21L port map( A => n2491, B => n1939, S => n2427, Z => n5725);
   U1294 : MUX21L port map( A => n2491, B => n868, S => n2428, Z => n5724);
   U1295 : MUX21L port map( A => n2491, B => n1938, S => n2429, Z => n5723);
   U1296 : MUX21L port map( A => n2491, B => n867, S => n2430, Z => n5722);
   U1297 : MUX21L port map( A => n1937, B => n2491, S => n2431, Z => n5721);
   U1298 : MUX21L port map( A => n866, B => n2491, S => n2432, Z => n5720);
   U1299 : MUX21L port map( A => n1936, B => n2491, S => n2433, Z => n5719);
   U1300 : MUX21L port map( A => n865, B => n2491, S => n2434, Z => n5718);
   U1301 : MUX21L port map( A => n2491, B => n1943, S => n2435, Z => n5717);
   U1302 : MUX21L port map( A => n2491, B => n872, S => n2436, Z => n5716);
   U1303 : MUX21L port map( A => n2491, B => n1942, S => n2437, Z => n5715);
   U1304 : MUX21L port map( A => n2491, B => n871, S => n2438, Z => n5714);
   U1305 : MUX21L port map( A => n1941, B => n2491, S => n2439, Z => n5713);
   U1306 : MUX21L port map( A => n870, B => n2491, S => n2440, Z => n5712);
   U1307 : MUX21L port map( A => n1940, B => n2491, S => n2441, Z => n5711);
   U1308 : MUX21L port map( A => n869, B => n2491, S => n2442, Z => n5710);
   U1309 : MUX21L port map( A => n2491, B => n1915, S => n2443, Z => n5709);
   U1310 : MUX21L port map( A => n2491, B => n844, S => n2444, Z => n5708);
   U1311 : MUX21L port map( A => n2491, B => n1914, S => n2445, Z => n5707);
   U1312 : MUX21L port map( A => n2491, B => n843, S => n2446, Z => n5706);
   U1313 : MUX21L port map( A => n1913, B => n2491, S => n2447, Z => n5705);
   U1314 : MUX21L port map( A => n842, B => n2491, S => n2448, Z => n5704);
   U1315 : MUX21L port map( A => n1912, B => n2491, S => n2449, Z => n5703);
   U1316 : MUX21L port map( A => n841, B => n2491, S => n2450, Z => n5702);
   U1317 : MUX21L port map( A => n2491, B => n1919, S => n2451, Z => n5701);
   U1318 : MUX21L port map( A => n2491, B => n848, S => n2452, Z => n5700);
   U1319 : MUX21L port map( A => n2491, B => n1918, S => n2453, Z => n5699);
   U1320 : MUX21L port map( A => n2491, B => n847, S => n2454, Z => n5698);
   U1321 : MUX21L port map( A => n1917, B => n2491, S => n2455, Z => n5697);
   U1322 : MUX21L port map( A => n846, B => n2491, S => n2456, Z => n5696);
   U1323 : MUX21L port map( A => n1916, B => n2491, S => n2457, Z => n5695);
   U1324 : MUX21L port map( A => n845, B => n2491, S => n2458, Z => n5694);
   U1325 : MUX21L port map( A => n2491, B => n1923, S => n2459, Z => n5693);
   U1326 : MUX21L port map( A => n2491, B => n852, S => n2460, Z => n5692);
   U1327 : MUX21L port map( A => n2491, B => n1922, S => n2461, Z => n5691);
   U1328 : MUX21L port map( A => n2491, B => n851, S => n2462, Z => n5690);
   U1329 : MUX21L port map( A => n1921, B => n2491, S => n2463, Z => n5689);
   U1330 : MUX21L port map( A => n850, B => n2491, S => n2464, Z => n5688);
   U1331 : MUX21L port map( A => n1920, B => n2491, S => n2465, Z => n5687);
   U1332 : MUX21L port map( A => n849, B => n2491, S => n2466, Z => n5686);
   U1333 : MUX21L port map( A => n2491, B => n1927, S => n2467, Z => n5685);
   U1334 : MUX21L port map( A => n2491, B => n856, S => n2468, Z => n5684);
   U1335 : MUX21L port map( A => n2491, B => n1926, S => n2469, Z => n5683);
   U1336 : MUX21L port map( A => n2491, B => n855, S => n2470, Z => n5682);
   U1337 : MUX21L port map( A => n1925, B => n2491, S => n2471, Z => n5681);
   U1338 : MUX21L port map( A => n854, B => n2491, S => n2472, Z => n5680);
   U1339 : MUX21L port map( A => n1924, B => n2491, S => n2473, Z => n5679);
   U1340 : MUX21L port map( A => n853, B => n2491, S => n2474, Z => n5678);
   U1341 : AO2 port map( A => v_TEMP_VECTOR_17_port, B => n2475, C => 
                           v_KEY32_IN_17_port, D => n2476, Z => n2491);
   U1342 : MUX21L port map( A => n2492, B => n2059, S => n2411, Z => n5677);
   U1343 : MUX21L port map( A => n2492, B => n988, S => n2412, Z => n5676);
   U1344 : MUX21L port map( A => n2492, B => n2058, S => n2413, Z => n5675);
   U1345 : MUX21L port map( A => n2492, B => n987, S => n2414, Z => n5674);
   U1346 : MUX21L port map( A => n2057, B => n2492, S => n2415, Z => n5673);
   U1347 : MUX21L port map( A => n986, B => n2492, S => n2416, Z => n5672);
   U1348 : MUX21L port map( A => n2056, B => n2492, S => n2417, Z => n5671);
   U1349 : MUX21L port map( A => n985, B => n2492, S => n2418, Z => n5670);
   U1350 : MUX21L port map( A => n2492, B => n2063, S => n2419, Z => n5669);
   U1351 : MUX21L port map( A => n2492, B => n992, S => n2420, Z => n5668);
   U1352 : MUX21L port map( A => n2492, B => n2062, S => n2421, Z => n5667);
   U1353 : MUX21L port map( A => n2492, B => n991, S => n2422, Z => n5666);
   U1354 : MUX21L port map( A => n2061, B => n2492, S => n2423, Z => n5665);
   U1355 : MUX21L port map( A => n990, B => n2492, S => n2424, Z => n5664);
   U1356 : MUX21L port map( A => n2060, B => n2492, S => n2425, Z => n5663);
   U1357 : MUX21L port map( A => n989, B => n2492, S => n2426, Z => n5662);
   U1358 : MUX21L port map( A => n2492, B => n2067, S => n2427, Z => n5661);
   U1359 : MUX21L port map( A => n2492, B => n996, S => n2428, Z => n5660);
   U1360 : MUX21L port map( A => n2492, B => n2066, S => n2429, Z => n5659);
   U1361 : MUX21L port map( A => n2492, B => n995, S => n2430, Z => n5658);
   U1362 : MUX21L port map( A => n2065, B => n2492, S => n2431, Z => n5657);
   U1363 : MUX21L port map( A => n994, B => n2492, S => n2432, Z => n5656);
   U1364 : MUX21L port map( A => n2064, B => n2492, S => n2433, Z => n5655);
   U1365 : MUX21L port map( A => n993, B => n2492, S => n2434, Z => n5654);
   U1366 : MUX21L port map( A => n2492, B => n2071, S => n2435, Z => n5653);
   U1367 : MUX21L port map( A => n2492, B => n1000, S => n2436, Z => n5652);
   U1368 : MUX21L port map( A => n2492, B => n2070, S => n2437, Z => n5651);
   U1369 : MUX21L port map( A => n2492, B => n999, S => n2438, Z => n5650);
   U1370 : MUX21L port map( A => n2069, B => n2492, S => n2439, Z => n5649);
   U1371 : MUX21L port map( A => n998, B => n2492, S => n2440, Z => n5648);
   U1372 : MUX21L port map( A => n2068, B => n2492, S => n2441, Z => n5647);
   U1373 : MUX21L port map( A => n997, B => n2492, S => n2442, Z => n5646);
   U1374 : MUX21L port map( A => n2492, B => n2043, S => n2443, Z => n5645);
   U1375 : MUX21L port map( A => n2492, B => n972, S => n2444, Z => n5644);
   U1376 : MUX21L port map( A => n2492, B => n2042, S => n2445, Z => n5643);
   U1377 : MUX21L port map( A => n2492, B => n971, S => n2446, Z => n5642);
   U1378 : MUX21L port map( A => n2041, B => n2492, S => n2447, Z => n5641);
   U1379 : MUX21L port map( A => n970, B => n2492, S => n2448, Z => n5640);
   U1380 : MUX21L port map( A => n2040, B => n2492, S => n2449, Z => n5639);
   U1381 : MUX21L port map( A => n969, B => n2492, S => n2450, Z => n5638);
   U1382 : MUX21L port map( A => n2492, B => n2047, S => n2451, Z => n5637);
   U1383 : MUX21L port map( A => n2492, B => n976, S => n2452, Z => n5636);
   U1384 : MUX21L port map( A => n2492, B => n2046, S => n2453, Z => n5635);
   U1385 : MUX21L port map( A => n2492, B => n975, S => n2454, Z => n5634);
   U1386 : MUX21L port map( A => n2045, B => n2492, S => n2455, Z => n5633);
   U1387 : MUX21L port map( A => n974, B => n2492, S => n2456, Z => n5632);
   U1388 : MUX21L port map( A => n2044, B => n2492, S => n2457, Z => n5631);
   U1389 : MUX21L port map( A => n973, B => n2492, S => n2458, Z => n5630);
   U1390 : MUX21L port map( A => n2492, B => n2051, S => n2459, Z => n5629);
   U1391 : MUX21L port map( A => n2492, B => n980, S => n2460, Z => n5628);
   U1392 : MUX21L port map( A => n2492, B => n2050, S => n2461, Z => n5627);
   U1393 : MUX21L port map( A => n2492, B => n979, S => n2462, Z => n5626);
   U1394 : MUX21L port map( A => n2049, B => n2492, S => n2463, Z => n5625);
   U1395 : MUX21L port map( A => n978, B => n2492, S => n2464, Z => n5624);
   U1396 : MUX21L port map( A => n2048, B => n2492, S => n2465, Z => n5623);
   U1397 : MUX21L port map( A => n977, B => n2492, S => n2466, Z => n5622);
   U1398 : MUX21L port map( A => n2492, B => n2055, S => n2467, Z => n5621);
   U1399 : MUX21L port map( A => n2492, B => n984, S => n2468, Z => n5620);
   U1400 : MUX21L port map( A => n2492, B => n2054, S => n2469, Z => n5619);
   U1401 : MUX21L port map( A => n2492, B => n983, S => n2470, Z => n5618);
   U1402 : MUX21L port map( A => n2053, B => n2492, S => n2471, Z => n5617);
   U1403 : MUX21L port map( A => n982, B => n2492, S => n2472, Z => n5616);
   U1404 : MUX21L port map( A => n2052, B => n2492, S => n2473, Z => n5615);
   U1405 : MUX21L port map( A => n981, B => n2492, S => n2474, Z => n5614);
   U1406 : AO2 port map( A => v_TEMP_VECTOR_16_port, B => n2475, C => 
                           v_KEY32_IN_16_port, D => n2476, Z => n2492);
   U1407 : MUX21L port map( A => n2493, B => n1195, S => n2411, Z => n5613);
   U1408 : MUX21L port map( A => n2493, B => n124, S => n2412, Z => n5612);
   U1409 : MUX21L port map( A => n2493, B => n1194, S => n2413, Z => n5611);
   U1410 : MUX21L port map( A => n2493, B => n123, S => n2414, Z => n5610);
   U1411 : MUX21L port map( A => n1193, B => n2493, S => n2415, Z => n5609);
   U1412 : MUX21L port map( A => n122, B => n2493, S => n2416, Z => n5608);
   U1413 : MUX21L port map( A => n1192, B => n2493, S => n2417, Z => n5607);
   U1414 : MUX21L port map( A => n121, B => n2493, S => n2418, Z => n5606);
   U1415 : MUX21L port map( A => n2493, B => n1199, S => n2419, Z => n5605);
   U1416 : MUX21L port map( A => n2493, B => n128, S => n2420, Z => n5604);
   U1417 : MUX21L port map( A => n2493, B => n1198, S => n2421, Z => n5603);
   U1418 : MUX21L port map( A => n2493, B => n127, S => n2422, Z => n5602);
   U1419 : MUX21L port map( A => n1197, B => n2493, S => n2423, Z => n5601);
   U1420 : MUX21L port map( A => n126, B => n2493, S => n2424, Z => n5600);
   U1421 : MUX21L port map( A => n1196, B => n2493, S => n2425, Z => n5599);
   U1422 : MUX21L port map( A => n125, B => n2493, S => n2426, Z => n5598);
   U1423 : MUX21L port map( A => n2493, B => n1203, S => n2427, Z => n5597);
   U1424 : MUX21L port map( A => n2493, B => n132, S => n2428, Z => n5596);
   U1425 : MUX21L port map( A => n2493, B => n1202, S => n2429, Z => n5595);
   U1426 : MUX21L port map( A => n2493, B => n131, S => n2430, Z => n5594);
   U1427 : MUX21L port map( A => n1201, B => n2493, S => n2431, Z => n5593);
   U1428 : MUX21L port map( A => n130, B => n2493, S => n2432, Z => n5592);
   U1429 : MUX21L port map( A => n1200, B => n2493, S => n2433, Z => n5591);
   U1430 : MUX21L port map( A => n129, B => n2493, S => n2434, Z => n5590);
   U1431 : MUX21L port map( A => n2493, B => n1207, S => n2435, Z => n5589);
   U1432 : MUX21L port map( A => n2493, B => n136, S => n2436, Z => n5588);
   U1433 : MUX21L port map( A => n2493, B => n1206, S => n2437, Z => n5587);
   U1434 : MUX21L port map( A => n2493, B => n135, S => n2438, Z => n5586);
   U1435 : MUX21L port map( A => n1205, B => n2493, S => n2439, Z => n5585);
   U1436 : MUX21L port map( A => n134, B => n2493, S => n2440, Z => n5584);
   U1437 : MUX21L port map( A => n1204, B => n2493, S => n2441, Z => n5583);
   U1438 : MUX21L port map( A => n133, B => n2493, S => n2442, Z => n5582);
   U1439 : MUX21L port map( A => n2493, B => n1179, S => n2443, Z => n5581);
   U1440 : MUX21L port map( A => n2493, B => n108, S => n2444, Z => n5580);
   U1441 : MUX21L port map( A => n2493, B => n1178, S => n2445, Z => n5579);
   U1442 : MUX21L port map( A => n2493, B => n107, S => n2446, Z => n5578);
   U1443 : MUX21L port map( A => n1177, B => n2493, S => n2447, Z => n5577);
   U1444 : MUX21L port map( A => n106, B => n2493, S => n2448, Z => n5576);
   U1445 : MUX21L port map( A => n1176, B => n2493, S => n2449, Z => n5575);
   U1446 : MUX21L port map( A => n105, B => n2493, S => n2450, Z => n5574);
   U1447 : MUX21L port map( A => n2493, B => n1183, S => n2451, Z => n5573);
   U1448 : MUX21L port map( A => n2493, B => n112, S => n2452, Z => n5572);
   U1449 : MUX21L port map( A => n2493, B => n1182, S => n2453, Z => n5571);
   U1450 : MUX21L port map( A => n2493, B => n111, S => n2454, Z => n5570);
   U1451 : MUX21L port map( A => n1181, B => n2493, S => n2455, Z => n5569);
   U1452 : MUX21L port map( A => n110, B => n2493, S => n2456, Z => n5568);
   U1453 : MUX21L port map( A => n1180, B => n2493, S => n2457, Z => n5567);
   U1454 : MUX21L port map( A => n109, B => n2493, S => n2458, Z => n5566);
   U1455 : MUX21L port map( A => n2493, B => n1187, S => n2459, Z => n5565);
   U1456 : MUX21L port map( A => n2493, B => n116, S => n2460, Z => n5564);
   U1457 : MUX21L port map( A => n2493, B => n1186, S => n2461, Z => n5563);
   U1458 : MUX21L port map( A => n2493, B => n115, S => n2462, Z => n5562);
   U1459 : MUX21L port map( A => n1185, B => n2493, S => n2463, Z => n5561);
   U1460 : MUX21L port map( A => n114, B => n2493, S => n2464, Z => n5560);
   U1461 : MUX21L port map( A => n1184, B => n2493, S => n2465, Z => n5559);
   U1462 : MUX21L port map( A => n113, B => n2493, S => n2466, Z => n5558);
   U1463 : MUX21L port map( A => n2493, B => n1191, S => n2467, Z => n5557);
   U1464 : MUX21L port map( A => n2493, B => n120, S => n2468, Z => n5556);
   U1465 : MUX21L port map( A => n2493, B => n1190, S => n2469, Z => n5555);
   U1466 : MUX21L port map( A => n2493, B => n119, S => n2470, Z => n5554);
   U1467 : MUX21L port map( A => n1189, B => n2493, S => n2471, Z => n5553);
   U1468 : MUX21L port map( A => n118, B => n2493, S => n2472, Z => n5552);
   U1469 : MUX21L port map( A => n1188, B => n2493, S => n2473, Z => n5551);
   U1470 : MUX21L port map( A => n117, B => n2493, S => n2474, Z => n5550);
   U1471 : AO2 port map( A => v_TEMP_VECTOR_15_port, B => n2475, C => 
                           v_KEY32_IN_15_port, D => n2476, Z => n2493);
   U1472 : MUX21L port map( A => n2494, B => n1323, S => n2411, Z => n5549);
   U1473 : MUX21L port map( A => n2494, B => n252, S => n2412, Z => n5548);
   U1474 : MUX21L port map( A => n2494, B => n1322, S => n2413, Z => n5547);
   U1475 : MUX21L port map( A => n2494, B => n251, S => n2414, Z => n5546);
   U1476 : MUX21L port map( A => n1321, B => n2494, S => n2415, Z => n5545);
   U1477 : MUX21L port map( A => n250, B => n2494, S => n2416, Z => n5544);
   U1478 : MUX21L port map( A => n1320, B => n2494, S => n2417, Z => n5543);
   U1479 : MUX21L port map( A => n249, B => n2494, S => n2418, Z => n5542);
   U1480 : MUX21L port map( A => n2494, B => n1327, S => n2419, Z => n5541);
   U1481 : MUX21L port map( A => n2494, B => n256, S => n2420, Z => n5540);
   U1482 : MUX21L port map( A => n2494, B => n1326, S => n2421, Z => n5539);
   U1483 : MUX21L port map( A => n2494, B => n255, S => n2422, Z => n5538);
   U1484 : MUX21L port map( A => n1325, B => n2494, S => n2423, Z => n5537);
   U1485 : MUX21L port map( A => n254, B => n2494, S => n2424, Z => n5536);
   U1486 : MUX21L port map( A => n1324, B => n2494, S => n2425, Z => n5535);
   U1487 : MUX21L port map( A => n253, B => n2494, S => n2426, Z => n5534);
   U1488 : MUX21L port map( A => n2494, B => n1331, S => n2427, Z => n5533);
   U1489 : MUX21L port map( A => n2494, B => n260, S => n2428, Z => n5532);
   U1490 : MUX21L port map( A => n2494, B => n1330, S => n2429, Z => n5531);
   U1491 : MUX21L port map( A => n2494, B => n259, S => n2430, Z => n5530);
   U1492 : MUX21L port map( A => n1329, B => n2494, S => n2431, Z => n5529);
   U1493 : MUX21L port map( A => n258, B => n2494, S => n2432, Z => n5528);
   U1494 : MUX21L port map( A => n1328, B => n2494, S => n2433, Z => n5527);
   U1495 : MUX21L port map( A => n257, B => n2494, S => n2434, Z => n5526);
   U1496 : MUX21L port map( A => n2494, B => n1335, S => n2435, Z => n5525);
   U1497 : MUX21L port map( A => n2494, B => n264, S => n2436, Z => n5524);
   U1498 : MUX21L port map( A => n2494, B => n1334, S => n2437, Z => n5523);
   U1499 : MUX21L port map( A => n2494, B => n263, S => n2438, Z => n5522);
   U1500 : MUX21L port map( A => n1333, B => n2494, S => n2439, Z => n5521);
   U1501 : MUX21L port map( A => n262, B => n2494, S => n2440, Z => n5520);
   U1502 : MUX21L port map( A => n1332, B => n2494, S => n2441, Z => n5519);
   U1503 : MUX21L port map( A => n261, B => n2494, S => n2442, Z => n5518);
   U1504 : MUX21L port map( A => n2494, B => n1307, S => n2443, Z => n5517);
   U1505 : MUX21L port map( A => n2494, B => n236, S => n2444, Z => n5516);
   U1506 : MUX21L port map( A => n2494, B => n1306, S => n2445, Z => n5515);
   U1507 : MUX21L port map( A => n2494, B => n235, S => n2446, Z => n5514);
   U1508 : MUX21L port map( A => n1305, B => n2494, S => n2447, Z => n5513);
   U1509 : MUX21L port map( A => n234, B => n2494, S => n2448, Z => n5512);
   U1510 : MUX21L port map( A => n1304, B => n2494, S => n2449, Z => n5511);
   U1511 : MUX21L port map( A => n233, B => n2494, S => n2450, Z => n5510);
   U1512 : MUX21L port map( A => n2494, B => n1311, S => n2451, Z => n5509);
   U1513 : MUX21L port map( A => n2494, B => n240, S => n2452, Z => n5508);
   U1514 : MUX21L port map( A => n2494, B => n1310, S => n2453, Z => n5507);
   U1515 : MUX21L port map( A => n2494, B => n239, S => n2454, Z => n5506);
   U1516 : MUX21L port map( A => n1309, B => n2494, S => n2455, Z => n5505);
   U1517 : MUX21L port map( A => n238, B => n2494, S => n2456, Z => n5504);
   U1518 : MUX21L port map( A => n1308, B => n2494, S => n2457, Z => n5503);
   U1519 : MUX21L port map( A => n237, B => n2494, S => n2458, Z => n5502);
   U1520 : MUX21L port map( A => n2494, B => n1315, S => n2459, Z => n5501);
   U1521 : MUX21L port map( A => n2494, B => n244, S => n2460, Z => n5500);
   U1522 : MUX21L port map( A => n2494, B => n1314, S => n2461, Z => n5499);
   U1523 : MUX21L port map( A => n2494, B => n243, S => n2462, Z => n5498);
   U1524 : MUX21L port map( A => n1313, B => n2494, S => n2463, Z => n5497);
   U1525 : MUX21L port map( A => n242, B => n2494, S => n2464, Z => n5496);
   U1526 : MUX21L port map( A => n1312, B => n2494, S => n2465, Z => n5495);
   U1527 : MUX21L port map( A => n241, B => n2494, S => n2466, Z => n5494);
   U1528 : MUX21L port map( A => n2494, B => n1319, S => n2467, Z => n5493);
   U1529 : MUX21L port map( A => n2494, B => n248, S => n2468, Z => n5492);
   U1530 : MUX21L port map( A => n2494, B => n1318, S => n2469, Z => n5491);
   U1531 : MUX21L port map( A => n2494, B => n247, S => n2470, Z => n5490);
   U1532 : MUX21L port map( A => n1317, B => n2494, S => n2471, Z => n5489);
   U1533 : MUX21L port map( A => n246, B => n2494, S => n2472, Z => n5488);
   U1534 : MUX21L port map( A => n1316, B => n2494, S => n2473, Z => n5487);
   U1535 : MUX21L port map( A => n245, B => n2494, S => n2474, Z => n5486);
   U1536 : AO2 port map( A => v_TEMP_VECTOR_14_port, B => n2475, C => 
                           v_KEY32_IN_14_port, D => n2476, Z => n2494);
   U1537 : MUX21L port map( A => n2495, B => n1451, S => n2411, Z => n5485);
   U1538 : MUX21L port map( A => n2495, B => n380, S => n2412, Z => n5484);
   U1539 : MUX21L port map( A => n2495, B => n1450, S => n2413, Z => n5483);
   U1540 : MUX21L port map( A => n2495, B => n379, S => n2414, Z => n5482);
   U1541 : MUX21L port map( A => n1449, B => n2495, S => n2415, Z => n5481);
   U1542 : MUX21L port map( A => n378, B => n2495, S => n2416, Z => n5480);
   U1543 : MUX21L port map( A => n1448, B => n2495, S => n2417, Z => n5479);
   U1544 : MUX21L port map( A => n377, B => n2495, S => n2418, Z => n5478);
   U1545 : MUX21L port map( A => n2495, B => n1455, S => n2419, Z => n5477);
   U1546 : MUX21L port map( A => n2495, B => n384, S => n2420, Z => n5476);
   U1547 : MUX21L port map( A => n2495, B => n1454, S => n2421, Z => n5475);
   U1548 : MUX21L port map( A => n2495, B => n383, S => n2422, Z => n5474);
   U1549 : MUX21L port map( A => n1453, B => n2495, S => n2423, Z => n5473);
   U1550 : MUX21L port map( A => n382, B => n2495, S => n2424, Z => n5472);
   U1551 : MUX21L port map( A => n1452, B => n2495, S => n2425, Z => n5471);
   U1552 : MUX21L port map( A => n381, B => n2495, S => n2426, Z => n5470);
   U1553 : MUX21L port map( A => n2495, B => n1459, S => n2427, Z => n5469);
   U1554 : MUX21L port map( A => n2495, B => n388, S => n2428, Z => n5468);
   U1555 : MUX21L port map( A => n2495, B => n1458, S => n2429, Z => n5467);
   U1556 : MUX21L port map( A => n2495, B => n387, S => n2430, Z => n5466);
   U1557 : MUX21L port map( A => n1457, B => n2495, S => n2431, Z => n5465);
   U1558 : MUX21L port map( A => n386, B => n2495, S => n2432, Z => n5464);
   U1559 : MUX21L port map( A => n1456, B => n2495, S => n2433, Z => n5463);
   U1560 : MUX21L port map( A => n385, B => n2495, S => n2434, Z => n5462);
   U1561 : MUX21L port map( A => n2495, B => n1463, S => n2435, Z => n5461);
   U1562 : MUX21L port map( A => n2495, B => n392, S => n2436, Z => n5460);
   U1563 : MUX21L port map( A => n2495, B => n1462, S => n2437, Z => n5459);
   U1564 : MUX21L port map( A => n2495, B => n391, S => n2438, Z => n5458);
   U1565 : MUX21L port map( A => n1461, B => n2495, S => n2439, Z => n5457);
   U1566 : MUX21L port map( A => n390, B => n2495, S => n2440, Z => n5456);
   U1567 : MUX21L port map( A => n1460, B => n2495, S => n2441, Z => n5455);
   U1568 : MUX21L port map( A => n389, B => n2495, S => n2442, Z => n5454);
   U1569 : MUX21L port map( A => n2495, B => n1435, S => n2443, Z => n5453);
   U1570 : MUX21L port map( A => n2495, B => n364, S => n2444, Z => n5452);
   U1571 : MUX21L port map( A => n2495, B => n1434, S => n2445, Z => n5451);
   U1572 : MUX21L port map( A => n2495, B => n363, S => n2446, Z => n5450);
   U1573 : MUX21L port map( A => n1433, B => n2495, S => n2447, Z => n5449);
   U1574 : MUX21L port map( A => n362, B => n2495, S => n2448, Z => n5448);
   U1575 : MUX21L port map( A => n1432, B => n2495, S => n2449, Z => n5447);
   U1576 : MUX21L port map( A => n361, B => n2495, S => n2450, Z => n5446);
   U1577 : MUX21L port map( A => n2495, B => n1439, S => n2451, Z => n5445);
   U1578 : MUX21L port map( A => n2495, B => n368, S => n2452, Z => n5444);
   U1579 : MUX21L port map( A => n2495, B => n1438, S => n2453, Z => n5443);
   U1580 : MUX21L port map( A => n2495, B => n367, S => n2454, Z => n5442);
   U1581 : MUX21L port map( A => n1437, B => n2495, S => n2455, Z => n5441);
   U1582 : MUX21L port map( A => n366, B => n2495, S => n2456, Z => n5440);
   U1583 : MUX21L port map( A => n1436, B => n2495, S => n2457, Z => n5439);
   U1584 : MUX21L port map( A => n365, B => n2495, S => n2458, Z => n5438);
   U1585 : MUX21L port map( A => n2495, B => n1443, S => n2459, Z => n5437);
   U1586 : MUX21L port map( A => n2495, B => n372, S => n2460, Z => n5436);
   U1587 : MUX21L port map( A => n2495, B => n1442, S => n2461, Z => n5435);
   U1588 : MUX21L port map( A => n2495, B => n371, S => n2462, Z => n5434);
   U1589 : MUX21L port map( A => n1441, B => n2495, S => n2463, Z => n5433);
   U1590 : MUX21L port map( A => n370, B => n2495, S => n2464, Z => n5432);
   U1591 : MUX21L port map( A => n1440, B => n2495, S => n2465, Z => n5431);
   U1592 : MUX21L port map( A => n369, B => n2495, S => n2466, Z => n5430);
   U1593 : MUX21L port map( A => n2495, B => n1447, S => n2467, Z => n5429);
   U1594 : MUX21L port map( A => n2495, B => n376, S => n2468, Z => n5428);
   U1595 : MUX21L port map( A => n2495, B => n1446, S => n2469, Z => n5427);
   U1596 : MUX21L port map( A => n2495, B => n375, S => n2470, Z => n5426);
   U1597 : MUX21L port map( A => n1445, B => n2495, S => n2471, Z => n5425);
   U1598 : MUX21L port map( A => n374, B => n2495, S => n2472, Z => n5424);
   U1599 : MUX21L port map( A => n1444, B => n2495, S => n2473, Z => n5423);
   U1600 : MUX21L port map( A => n373, B => n2495, S => n2474, Z => n5422);
   U1601 : AO2 port map( A => v_TEMP_VECTOR_13_port, B => n2475, C => 
                           v_KEY32_IN_13_port, D => n2476, Z => n2495);
   U1602 : MUX21L port map( A => n2496, B => n1579, S => n2411, Z => n5421);
   U1603 : MUX21L port map( A => n2496, B => n508, S => n2412, Z => n5420);
   U1604 : MUX21L port map( A => n2496, B => n1578, S => n2413, Z => n5419);
   U1605 : MUX21L port map( A => n2496, B => n507, S => n2414, Z => n5418);
   U1606 : MUX21L port map( A => n1577, B => n2496, S => n2415, Z => n5417);
   U1607 : MUX21L port map( A => n506, B => n2496, S => n2416, Z => n5416);
   U1608 : MUX21L port map( A => n1576, B => n2496, S => n2417, Z => n5415);
   U1609 : MUX21L port map( A => n505, B => n2496, S => n2418, Z => n5414);
   U1610 : MUX21L port map( A => n2496, B => n1583, S => n2419, Z => n5413);
   U1611 : MUX21L port map( A => n2496, B => n512, S => n2420, Z => n5412);
   U1612 : MUX21L port map( A => n2496, B => n1582, S => n2421, Z => n5411);
   U1613 : MUX21L port map( A => n2496, B => n511, S => n2422, Z => n5410);
   U1614 : MUX21L port map( A => n1581, B => n2496, S => n2423, Z => n5409);
   U1615 : MUX21L port map( A => n510, B => n2496, S => n2424, Z => n5408);
   U1616 : MUX21L port map( A => n1580, B => n2496, S => n2425, Z => n5407);
   U1617 : MUX21L port map( A => n509, B => n2496, S => n2426, Z => n5406);
   U1618 : MUX21L port map( A => n2496, B => n1587, S => n2427, Z => n5405);
   U1619 : MUX21L port map( A => n2496, B => n516, S => n2428, Z => n5404);
   U1620 : MUX21L port map( A => n2496, B => n1586, S => n2429, Z => n5403);
   U1621 : MUX21L port map( A => n2496, B => n515, S => n2430, Z => n5402);
   U1622 : MUX21L port map( A => n1585, B => n2496, S => n2431, Z => n5401);
   U1623 : MUX21L port map( A => n514, B => n2496, S => n2432, Z => n5400);
   U1624 : MUX21L port map( A => n1584, B => n2496, S => n2433, Z => n5399);
   U1625 : MUX21L port map( A => n513, B => n2496, S => n2434, Z => n5398);
   U1626 : MUX21L port map( A => n2496, B => n1591, S => n2435, Z => n5397);
   U1627 : MUX21L port map( A => n2496, B => n520, S => n2436, Z => n5396);
   U1628 : MUX21L port map( A => n2496, B => n1590, S => n2437, Z => n5395);
   U1629 : MUX21L port map( A => n2496, B => n519, S => n2438, Z => n5394);
   U1630 : MUX21L port map( A => n1589, B => n2496, S => n2439, Z => n5393);
   U1631 : MUX21L port map( A => n518, B => n2496, S => n2440, Z => n5392);
   U1632 : MUX21L port map( A => n1588, B => n2496, S => n2441, Z => n5391);
   U1633 : MUX21L port map( A => n517, B => n2496, S => n2442, Z => n5390);
   U1634 : MUX21L port map( A => n2496, B => n1563, S => n2443, Z => n5389);
   U1635 : MUX21L port map( A => n2496, B => n492, S => n2444, Z => n5388);
   U1636 : MUX21L port map( A => n2496, B => n1562, S => n2445, Z => n5387);
   U1637 : MUX21L port map( A => n2496, B => n491, S => n2446, Z => n5386);
   U1638 : MUX21L port map( A => n1561, B => n2496, S => n2447, Z => n5385);
   U1639 : MUX21L port map( A => n490, B => n2496, S => n2448, Z => n5384);
   U1640 : MUX21L port map( A => n1560, B => n2496, S => n2449, Z => n5383);
   U1641 : MUX21L port map( A => n489, B => n2496, S => n2450, Z => n5382);
   U1642 : MUX21L port map( A => n2496, B => n1567, S => n2451, Z => n5381);
   U1643 : MUX21L port map( A => n2496, B => n496, S => n2452, Z => n5380);
   U1644 : MUX21L port map( A => n2496, B => n1566, S => n2453, Z => n5379);
   U1645 : MUX21L port map( A => n2496, B => n495, S => n2454, Z => n5378);
   U1646 : MUX21L port map( A => n1565, B => n2496, S => n2455, Z => n5377);
   U1647 : MUX21L port map( A => n494, B => n2496, S => n2456, Z => n5376);
   U1648 : MUX21L port map( A => n1564, B => n2496, S => n2457, Z => n5375);
   U1649 : MUX21L port map( A => n493, B => n2496, S => n2458, Z => n5374);
   U1650 : MUX21L port map( A => n2496, B => n1571, S => n2459, Z => n5373);
   U1651 : MUX21L port map( A => n2496, B => n500, S => n2460, Z => n5372);
   U1652 : MUX21L port map( A => n2496, B => n1570, S => n2461, Z => n5371);
   U1653 : MUX21L port map( A => n2496, B => n499, S => n2462, Z => n5370);
   U1654 : MUX21L port map( A => n1569, B => n2496, S => n2463, Z => n5369);
   U1655 : MUX21L port map( A => n498, B => n2496, S => n2464, Z => n5368);
   U1656 : MUX21L port map( A => n1568, B => n2496, S => n2465, Z => n5367);
   U1657 : MUX21L port map( A => n497, B => n2496, S => n2466, Z => n5366);
   U1658 : MUX21L port map( A => n2496, B => n1575, S => n2467, Z => n5365);
   U1659 : MUX21L port map( A => n2496, B => n504, S => n2468, Z => n5364);
   U1660 : MUX21L port map( A => n2496, B => n1574, S => n2469, Z => n5363);
   U1661 : MUX21L port map( A => n2496, B => n503, S => n2470, Z => n5362);
   U1662 : MUX21L port map( A => n1573, B => n2496, S => n2471, Z => n5361);
   U1663 : MUX21L port map( A => n502, B => n2496, S => n2472, Z => n5360);
   U1664 : MUX21L port map( A => n1572, B => n2496, S => n2473, Z => n5359);
   U1665 : MUX21L port map( A => n501, B => n2496, S => n2474, Z => n5358);
   U1666 : AO2 port map( A => v_TEMP_VECTOR_12_port, B => n2475, C => 
                           v_KEY32_IN_12_port, D => n2476, Z => n2496);
   U1667 : MUX21L port map( A => n2497, B => n1707, S => n2411, Z => n5357);
   U1668 : MUX21L port map( A => n2497, B => n636, S => n2412, Z => n5356);
   U1669 : MUX21L port map( A => n2497, B => n1706, S => n2413, Z => n5355);
   U1670 : MUX21L port map( A => n2497, B => n635, S => n2414, Z => n5354);
   U1671 : MUX21L port map( A => n1705, B => n2497, S => n2415, Z => n5353);
   U1672 : MUX21L port map( A => n634, B => n2497, S => n2416, Z => n5352);
   U1673 : MUX21L port map( A => n1704, B => n2497, S => n2417, Z => n5351);
   U1674 : MUX21L port map( A => n633, B => n2497, S => n2418, Z => n5350);
   U1675 : MUX21L port map( A => n2497, B => n1711, S => n2419, Z => n5349);
   U1676 : MUX21L port map( A => n2497, B => n640, S => n2420, Z => n5348);
   U1677 : MUX21L port map( A => n2497, B => n1710, S => n2421, Z => n5347);
   U1678 : MUX21L port map( A => n2497, B => n639, S => n2422, Z => n5346);
   U1679 : MUX21L port map( A => n1709, B => n2497, S => n2423, Z => n5345);
   U1680 : MUX21L port map( A => n638, B => n2497, S => n2424, Z => n5344);
   U1681 : MUX21L port map( A => n1708, B => n2497, S => n2425, Z => n5343);
   U1682 : MUX21L port map( A => n637, B => n2497, S => n2426, Z => n5342);
   U1683 : MUX21L port map( A => n2497, B => n1715, S => n2427, Z => n5341);
   U1684 : MUX21L port map( A => n2497, B => n644, S => n2428, Z => n5340);
   U1685 : MUX21L port map( A => n2497, B => n1714, S => n2429, Z => n5339);
   U1686 : MUX21L port map( A => n2497, B => n643, S => n2430, Z => n5338);
   U1687 : MUX21L port map( A => n1713, B => n2497, S => n2431, Z => n5337);
   U1688 : MUX21L port map( A => n642, B => n2497, S => n2432, Z => n5336);
   U1689 : MUX21L port map( A => n1712, B => n2497, S => n2433, Z => n5335);
   U1690 : MUX21L port map( A => n641, B => n2497, S => n2434, Z => n5334);
   U1691 : MUX21L port map( A => n2497, B => n1719, S => n2435, Z => n5333);
   U1692 : MUX21L port map( A => n2497, B => n648, S => n2436, Z => n5332);
   U1693 : MUX21L port map( A => n2497, B => n1718, S => n2437, Z => n5331);
   U1694 : MUX21L port map( A => n2497, B => n647, S => n2438, Z => n5330);
   U1695 : MUX21L port map( A => n1717, B => n2497, S => n2439, Z => n5329);
   U1696 : MUX21L port map( A => n646, B => n2497, S => n2440, Z => n5328);
   U1697 : MUX21L port map( A => n1716, B => n2497, S => n2441, Z => n5327);
   U1698 : MUX21L port map( A => n645, B => n2497, S => n2442, Z => n5326);
   U1699 : MUX21L port map( A => n2497, B => n1691, S => n2443, Z => n5325);
   U1700 : MUX21L port map( A => n2497, B => n620, S => n2444, Z => n5324);
   U1701 : MUX21L port map( A => n2497, B => n1690, S => n2445, Z => n5323);
   U1702 : MUX21L port map( A => n2497, B => n619, S => n2446, Z => n5322);
   U1703 : MUX21L port map( A => n1689, B => n2497, S => n2447, Z => n5321);
   U1704 : MUX21L port map( A => n618, B => n2497, S => n2448, Z => n5320);
   U1705 : MUX21L port map( A => n1688, B => n2497, S => n2449, Z => n5319);
   U1706 : MUX21L port map( A => n617, B => n2497, S => n2450, Z => n5318);
   U1707 : MUX21L port map( A => n2497, B => n1695, S => n2451, Z => n5317);
   U1708 : MUX21L port map( A => n2497, B => n624, S => n2452, Z => n5316);
   U1709 : MUX21L port map( A => n2497, B => n1694, S => n2453, Z => n5315);
   U1710 : MUX21L port map( A => n2497, B => n623, S => n2454, Z => n5314);
   U1711 : MUX21L port map( A => n1693, B => n2497, S => n2455, Z => n5313);
   U1712 : MUX21L port map( A => n622, B => n2497, S => n2456, Z => n5312);
   U1713 : MUX21L port map( A => n1692, B => n2497, S => n2457, Z => n5311);
   U1714 : MUX21L port map( A => n621, B => n2497, S => n2458, Z => n5310);
   U1715 : MUX21L port map( A => n2497, B => n1699, S => n2459, Z => n5309);
   U1716 : MUX21L port map( A => n2497, B => n628, S => n2460, Z => n5308);
   U1717 : MUX21L port map( A => n2497, B => n1698, S => n2461, Z => n5307);
   U1718 : MUX21L port map( A => n2497, B => n627, S => n2462, Z => n5306);
   U1719 : MUX21L port map( A => n1697, B => n2497, S => n2463, Z => n5305);
   U1720 : MUX21L port map( A => n626, B => n2497, S => n2464, Z => n5304);
   U1721 : MUX21L port map( A => n1696, B => n2497, S => n2465, Z => n5303);
   U1722 : MUX21L port map( A => n625, B => n2497, S => n2466, Z => n5302);
   U1723 : MUX21L port map( A => n2497, B => n1703, S => n2467, Z => n5301);
   U1724 : MUX21L port map( A => n2497, B => n632, S => n2468, Z => n5300);
   U1725 : MUX21L port map( A => n2497, B => n1702, S => n2469, Z => n5299);
   U1726 : MUX21L port map( A => n2497, B => n631, S => n2470, Z => n5298);
   U1727 : MUX21L port map( A => n1701, B => n2497, S => n2471, Z => n5297);
   U1728 : MUX21L port map( A => n630, B => n2497, S => n2472, Z => n5296);
   U1729 : MUX21L port map( A => n1700, B => n2497, S => n2473, Z => n5295);
   U1730 : MUX21L port map( A => n629, B => n2497, S => n2474, Z => n5294);
   U1731 : AO2 port map( A => v_TEMP_VECTOR_11_port, B => n2475, C => 
                           v_KEY32_IN_11_port, D => n2476, Z => n2497);
   U1732 : MUX21L port map( A => n2498, B => n1835, S => n2411, Z => n5293);
   U1733 : MUX21L port map( A => n2498, B => n764, S => n2412, Z => n5292);
   U1734 : MUX21L port map( A => n2498, B => n1834, S => n2413, Z => n5291);
   U1735 : MUX21L port map( A => n2498, B => n763, S => n2414, Z => n5290);
   U1736 : MUX21L port map( A => n1833, B => n2498, S => n2415, Z => n5289);
   U1737 : MUX21L port map( A => n762, B => n2498, S => n2416, Z => n5288);
   U1738 : MUX21L port map( A => n1832, B => n2498, S => n2417, Z => n5287);
   U1739 : MUX21L port map( A => n761, B => n2498, S => n2418, Z => n5286);
   U1740 : MUX21L port map( A => n2498, B => n1839, S => n2419, Z => n5285);
   U1741 : MUX21L port map( A => n2498, B => n768, S => n2420, Z => n5284);
   U1742 : MUX21L port map( A => n2498, B => n1838, S => n2421, Z => n5283);
   U1743 : MUX21L port map( A => n2498, B => n767, S => n2422, Z => n5282);
   U1744 : MUX21L port map( A => n1837, B => n2498, S => n2423, Z => n5281);
   U1745 : MUX21L port map( A => n766, B => n2498, S => n2424, Z => n5280);
   U1746 : MUX21L port map( A => n1836, B => n2498, S => n2425, Z => n5279);
   U1747 : MUX21L port map( A => n765, B => n2498, S => n2426, Z => n5278);
   U1748 : MUX21L port map( A => n2498, B => n1843, S => n2427, Z => n5277);
   U1749 : MUX21L port map( A => n2498, B => n772, S => n2428, Z => n5276);
   U1750 : MUX21L port map( A => n2498, B => n1842, S => n2429, Z => n5275);
   U1751 : MUX21L port map( A => n2498, B => n771, S => n2430, Z => n5274);
   U1752 : MUX21L port map( A => n1841, B => n2498, S => n2431, Z => n5273);
   U1753 : MUX21L port map( A => n770, B => n2498, S => n2432, Z => n5272);
   U1754 : MUX21L port map( A => n1840, B => n2498, S => n2433, Z => n5271);
   U1755 : MUX21L port map( A => n769, B => n2498, S => n2434, Z => n5270);
   U1756 : MUX21L port map( A => n2498, B => n1847, S => n2435, Z => n5269);
   U1757 : MUX21L port map( A => n2498, B => n776, S => n2436, Z => n5268);
   U1758 : MUX21L port map( A => n2498, B => n1846, S => n2437, Z => n5267);
   U1759 : MUX21L port map( A => n2498, B => n775, S => n2438, Z => n5266);
   U1760 : MUX21L port map( A => n1845, B => n2498, S => n2439, Z => n5265);
   U1761 : MUX21L port map( A => n774, B => n2498, S => n2440, Z => n5264);
   U1762 : MUX21L port map( A => n1844, B => n2498, S => n2441, Z => n5263);
   U1763 : MUX21L port map( A => n773, B => n2498, S => n2442, Z => n5262);
   U1764 : MUX21L port map( A => n2498, B => n1819, S => n2443, Z => n5261);
   U1765 : MUX21L port map( A => n2498, B => n748, S => n2444, Z => n5260);
   U1766 : MUX21L port map( A => n2498, B => n1818, S => n2445, Z => n5259);
   U1767 : MUX21L port map( A => n2498, B => n747, S => n2446, Z => n5258);
   U1768 : MUX21L port map( A => n1817, B => n2498, S => n2447, Z => n5257);
   U1769 : MUX21L port map( A => n746, B => n2498, S => n2448, Z => n5256);
   U1770 : MUX21L port map( A => n1816, B => n2498, S => n2449, Z => n5255);
   U1771 : MUX21L port map( A => n745, B => n2498, S => n2450, Z => n5254);
   U1772 : MUX21L port map( A => n2498, B => n1823, S => n2451, Z => n5253);
   U1773 : MUX21L port map( A => n2498, B => n752, S => n2452, Z => n5252);
   U1774 : MUX21L port map( A => n2498, B => n1822, S => n2453, Z => n5251);
   U1775 : MUX21L port map( A => n2498, B => n751, S => n2454, Z => n5250);
   U1776 : MUX21L port map( A => n1821, B => n2498, S => n2455, Z => n5249);
   U1777 : MUX21L port map( A => n750, B => n2498, S => n2456, Z => n5248);
   U1778 : MUX21L port map( A => n1820, B => n2498, S => n2457, Z => n5247);
   U1779 : MUX21L port map( A => n749, B => n2498, S => n2458, Z => n5246);
   U1780 : MUX21L port map( A => n2498, B => n1827, S => n2459, Z => n5245);
   U1781 : MUX21L port map( A => n2498, B => n756, S => n2460, Z => n5244);
   U1782 : MUX21L port map( A => n2498, B => n1826, S => n2461, Z => n5243);
   U1783 : MUX21L port map( A => n2498, B => n755, S => n2462, Z => n5242);
   U1784 : MUX21L port map( A => n1825, B => n2498, S => n2463, Z => n5241);
   U1785 : MUX21L port map( A => n754, B => n2498, S => n2464, Z => n5240);
   U1786 : MUX21L port map( A => n1824, B => n2498, S => n2465, Z => n5239);
   U1787 : MUX21L port map( A => n753, B => n2498, S => n2466, Z => n5238);
   U1788 : MUX21L port map( A => n2498, B => n1831, S => n2467, Z => n5237);
   U1789 : MUX21L port map( A => n2498, B => n760, S => n2468, Z => n5236);
   U1790 : MUX21L port map( A => n2498, B => n1830, S => n2469, Z => n5235);
   U1791 : MUX21L port map( A => n2498, B => n759, S => n2470, Z => n5234);
   U1792 : MUX21L port map( A => n1829, B => n2498, S => n2471, Z => n5233);
   U1793 : MUX21L port map( A => n758, B => n2498, S => n2472, Z => n5232);
   U1794 : MUX21L port map( A => n1828, B => n2498, S => n2473, Z => n5231);
   U1795 : MUX21L port map( A => n757, B => n2498, S => n2474, Z => n5230);
   U1796 : AO2 port map( A => v_TEMP_VECTOR_10_port, B => n2475, C => 
                           v_KEY32_IN_10_port, D => n2476, Z => n2498);
   U1797 : MUX21L port map( A => n2499, B => n1963, S => n2411, Z => n5229);
   U1798 : MUX21L port map( A => n2499, B => n892, S => n2412, Z => n5228);
   U1799 : MUX21L port map( A => n2499, B => n1962, S => n2413, Z => n5227);
   U1800 : MUX21L port map( A => n2499, B => n891, S => n2414, Z => n5226);
   U1801 : MUX21L port map( A => n1961, B => n2499, S => n2415, Z => n5225);
   U1802 : MUX21L port map( A => n890, B => n2499, S => n2416, Z => n5224);
   U1803 : MUX21L port map( A => n1960, B => n2499, S => n2417, Z => n5223);
   U1804 : MUX21L port map( A => n889, B => n2499, S => n2418, Z => n5222);
   U1805 : MUX21L port map( A => n2499, B => n1967, S => n2419, Z => n5221);
   U1806 : MUX21L port map( A => n2499, B => n896, S => n2420, Z => n5220);
   U1807 : MUX21L port map( A => n2499, B => n1966, S => n2421, Z => n5219);
   U1808 : MUX21L port map( A => n2499, B => n895, S => n2422, Z => n5218);
   U1809 : MUX21L port map( A => n1965, B => n2499, S => n2423, Z => n5217);
   U1810 : MUX21L port map( A => n894, B => n2499, S => n2424, Z => n5216);
   U1811 : MUX21L port map( A => n1964, B => n2499, S => n2425, Z => n5215);
   U1812 : MUX21L port map( A => n893, B => n2499, S => n2426, Z => n5214);
   U1813 : MUX21L port map( A => n2499, B => n1971, S => n2427, Z => n5213);
   U1814 : MUX21L port map( A => n2499, B => n900, S => n2428, Z => n5212);
   U1815 : MUX21L port map( A => n2499, B => n1970, S => n2429, Z => n5211);
   U1816 : MUX21L port map( A => n2499, B => n899, S => n2430, Z => n5210);
   U1817 : MUX21L port map( A => n1969, B => n2499, S => n2431, Z => n5209);
   U1818 : MUX21L port map( A => n898, B => n2499, S => n2432, Z => n5208);
   U1819 : MUX21L port map( A => n1968, B => n2499, S => n2433, Z => n5207);
   U1820 : MUX21L port map( A => n897, B => n2499, S => n2434, Z => n5206);
   U1821 : MUX21L port map( A => n2499, B => n1975, S => n2435, Z => n5205);
   U1822 : MUX21L port map( A => n2499, B => n904, S => n2436, Z => n5204);
   U1823 : MUX21L port map( A => n2499, B => n1974, S => n2437, Z => n5203);
   U1824 : MUX21L port map( A => n2499, B => n903, S => n2438, Z => n5202);
   U1825 : MUX21L port map( A => n1973, B => n2499, S => n2439, Z => n5201);
   U1826 : MUX21L port map( A => n902, B => n2499, S => n2440, Z => n5200);
   U1827 : MUX21L port map( A => n1972, B => n2499, S => n2441, Z => n5199);
   U1828 : MUX21L port map( A => n901, B => n2499, S => n2442, Z => n5198);
   U1829 : MUX21L port map( A => n2499, B => n1947, S => n2443, Z => n5197);
   U1830 : MUX21L port map( A => n2499, B => n876, S => n2444, Z => n5196);
   U1831 : MUX21L port map( A => n2499, B => n1946, S => n2445, Z => n5195);
   U1832 : MUX21L port map( A => n2499, B => n875, S => n2446, Z => n5194);
   U1833 : MUX21L port map( A => n1945, B => n2499, S => n2447, Z => n5193);
   U1834 : MUX21L port map( A => n874, B => n2499, S => n2448, Z => n5192);
   U1835 : MUX21L port map( A => n1944, B => n2499, S => n2449, Z => n5191);
   U1836 : MUX21L port map( A => n873, B => n2499, S => n2450, Z => n5190);
   U1837 : MUX21L port map( A => n2499, B => n1951, S => n2451, Z => n5189);
   U1838 : MUX21L port map( A => n2499, B => n880, S => n2452, Z => n5188);
   U1839 : MUX21L port map( A => n2499, B => n1950, S => n2453, Z => n5187);
   U1840 : MUX21L port map( A => n2499, B => n879, S => n2454, Z => n5186);
   U1841 : MUX21L port map( A => n1949, B => n2499, S => n2455, Z => n5185);
   U1842 : MUX21L port map( A => n878, B => n2499, S => n2456, Z => n5184);
   U1843 : MUX21L port map( A => n1948, B => n2499, S => n2457, Z => n5183);
   U1844 : MUX21L port map( A => n877, B => n2499, S => n2458, Z => n5182);
   U1845 : MUX21L port map( A => n2499, B => n1955, S => n2459, Z => n5181);
   U1846 : MUX21L port map( A => n2499, B => n884, S => n2460, Z => n5180);
   U1847 : MUX21L port map( A => n2499, B => n1954, S => n2461, Z => n5179);
   U1848 : MUX21L port map( A => n2499, B => n883, S => n2462, Z => n5178);
   U1849 : MUX21L port map( A => n1953, B => n2499, S => n2463, Z => n5177);
   U1850 : MUX21L port map( A => n882, B => n2499, S => n2464, Z => n5176);
   U1851 : MUX21L port map( A => n1952, B => n2499, S => n2465, Z => n5175);
   U1852 : MUX21L port map( A => n881, B => n2499, S => n2466, Z => n5174);
   U1853 : MUX21L port map( A => n2499, B => n1959, S => n2467, Z => n5173);
   U1854 : MUX21L port map( A => n2499, B => n888, S => n2468, Z => n5172);
   U1855 : MUX21L port map( A => n2499, B => n1958, S => n2469, Z => n5171);
   U1856 : MUX21L port map( A => n2499, B => n887, S => n2470, Z => n5170);
   U1857 : MUX21L port map( A => n1957, B => n2499, S => n2471, Z => n5169);
   U1858 : MUX21L port map( A => n886, B => n2499, S => n2472, Z => n5168);
   U1859 : MUX21L port map( A => n1956, B => n2499, S => n2473, Z => n5167);
   U1860 : MUX21L port map( A => n885, B => n2499, S => n2474, Z => n5166);
   U1861 : AO2 port map( A => v_TEMP_VECTOR_9_port, B => n2475, C => 
                           v_KEY32_IN_9_port, D => n2476, Z => n2499);
   U1862 : MUX21L port map( A => n2500, B => n2091, S => n2411, Z => n5165);
   U1863 : MUX21L port map( A => n2500, B => n1020, S => n2412, Z => n5164);
   U1864 : MUX21L port map( A => n2500, B => n2090, S => n2413, Z => n5163);
   U1865 : MUX21L port map( A => n2500, B => n1019, S => n2414, Z => n5162);
   U1866 : MUX21L port map( A => n2089, B => n2500, S => n2415, Z => n5161);
   U1867 : MUX21L port map( A => n1018, B => n2500, S => n2416, Z => n5160);
   U1868 : MUX21L port map( A => n2088, B => n2500, S => n2417, Z => n5159);
   U1869 : MUX21L port map( A => n1017, B => n2500, S => n2418, Z => n5158);
   U1870 : MUX21L port map( A => n2500, B => n2095, S => n2419, Z => n5157);
   U1871 : MUX21L port map( A => n2500, B => n1024, S => n2420, Z => n5156);
   U1872 : MUX21L port map( A => n2500, B => n2094, S => n2421, Z => n5155);
   U1873 : MUX21L port map( A => n2500, B => n1023, S => n2422, Z => n5154);
   U1874 : MUX21L port map( A => n2093, B => n2500, S => n2423, Z => n5153);
   U1875 : MUX21L port map( A => n1022, B => n2500, S => n2424, Z => n5152);
   U1876 : MUX21L port map( A => n2092, B => n2500, S => n2425, Z => n5151);
   U1877 : MUX21L port map( A => n1021, B => n2500, S => n2426, Z => n5150);
   U1878 : MUX21L port map( A => n2500, B => n2099, S => n2427, Z => n5149);
   U1879 : MUX21L port map( A => n2500, B => n1028, S => n2428, Z => n5148);
   U1880 : MUX21L port map( A => n2500, B => n2098, S => n2429, Z => n5147);
   U1881 : MUX21L port map( A => n2500, B => n1027, S => n2430, Z => n5146);
   U1882 : MUX21L port map( A => n2097, B => n2500, S => n2431, Z => n5145);
   U1883 : MUX21L port map( A => n1026, B => n2500, S => n2432, Z => n5144);
   U1884 : MUX21L port map( A => n2096, B => n2500, S => n2433, Z => n5143);
   U1885 : MUX21L port map( A => n1025, B => n2500, S => n2434, Z => n5142);
   U1886 : MUX21L port map( A => n2500, B => n2103, S => n2435, Z => n5141);
   U1887 : MUX21L port map( A => n2500, B => n1032, S => n2436, Z => n5140);
   U1888 : MUX21L port map( A => n2500, B => n2102, S => n2437, Z => n5139);
   U1889 : MUX21L port map( A => n2500, B => n1031, S => n2438, Z => n5138);
   U1890 : MUX21L port map( A => n2101, B => n2500, S => n2439, Z => n5137);
   U1891 : MUX21L port map( A => n1030, B => n2500, S => n2440, Z => n5136);
   U1892 : MUX21L port map( A => n2100, B => n2500, S => n2441, Z => n5135);
   U1893 : MUX21L port map( A => n1029, B => n2500, S => n2442, Z => n5134);
   U1894 : MUX21L port map( A => n2500, B => n2075, S => n2443, Z => n5133);
   U1895 : MUX21L port map( A => n2500, B => n1004, S => n2444, Z => n5132);
   U1896 : MUX21L port map( A => n2500, B => n2074, S => n2445, Z => n5131);
   U1897 : MUX21L port map( A => n2500, B => n1003, S => n2446, Z => n5130);
   U1898 : MUX21L port map( A => n2073, B => n2500, S => n2447, Z => n5129);
   U1899 : MUX21L port map( A => n1002, B => n2500, S => n2448, Z => n5128);
   U1900 : MUX21L port map( A => n2072, B => n2500, S => n2449, Z => n5127);
   U1901 : MUX21L port map( A => n1001, B => n2500, S => n2450, Z => n5126);
   U1902 : MUX21L port map( A => n2500, B => n2079, S => n2451, Z => n5125);
   U1903 : MUX21L port map( A => n2500, B => n1008, S => n2452, Z => n5124);
   U1904 : MUX21L port map( A => n2500, B => n2078, S => n2453, Z => n5123);
   U1905 : MUX21L port map( A => n2500, B => n1007, S => n2454, Z => n5122);
   U1906 : MUX21L port map( A => n2077, B => n2500, S => n2455, Z => n5121);
   U1907 : MUX21L port map( A => n1006, B => n2500, S => n2456, Z => n5120);
   U1908 : MUX21L port map( A => n2076, B => n2500, S => n2457, Z => n5119);
   U1909 : MUX21L port map( A => n1005, B => n2500, S => n2458, Z => n5118);
   U1910 : MUX21L port map( A => n2500, B => n2083, S => n2459, Z => n5117);
   U1911 : MUX21L port map( A => n2500, B => n1012, S => n2460, Z => n5116);
   U1912 : MUX21L port map( A => n2500, B => n2082, S => n2461, Z => n5115);
   U1913 : MUX21L port map( A => n2500, B => n1011, S => n2462, Z => n5114);
   U1914 : MUX21L port map( A => n2081, B => n2500, S => n2463, Z => n5113);
   U1915 : MUX21L port map( A => n1010, B => n2500, S => n2464, Z => n5112);
   U1916 : MUX21L port map( A => n2080, B => n2500, S => n2465, Z => n5111);
   U1917 : MUX21L port map( A => n1009, B => n2500, S => n2466, Z => n5110);
   U1918 : MUX21L port map( A => n2500, B => n2087, S => n2467, Z => n5109);
   U1919 : MUX21L port map( A => n2500, B => n1016, S => n2468, Z => n5108);
   U1920 : MUX21L port map( A => n2500, B => n2086, S => n2469, Z => n5107);
   U1921 : MUX21L port map( A => n2500, B => n1015, S => n2470, Z => n5106);
   U1922 : MUX21L port map( A => n2085, B => n2500, S => n2471, Z => n5105);
   U1923 : MUX21L port map( A => n1014, B => n2500, S => n2472, Z => n5104);
   U1924 : MUX21L port map( A => n2084, B => n2500, S => n2473, Z => n5103);
   U1925 : MUX21L port map( A => n1013, B => n2500, S => n2474, Z => n5102);
   U1926 : AO2 port map( A => v_TEMP_VECTOR_8_port, B => n2475, C => 
                           v_KEY32_IN_8_port, D => n2476, Z => n2500);
   U1927 : MUX21L port map( A => n2501, B => n1099, S => n2411, Z => n5101);
   U1928 : MUX21L port map( A => n2501, B => n28, S => n2412, Z => n5100);
   U1929 : MUX21L port map( A => n2501, B => n1098, S => n2413, Z => n5099);
   U1930 : MUX21L port map( A => n2501, B => n27, S => n2414, Z => n5098);
   U1931 : MUX21L port map( A => n1097, B => n2501, S => n2415, Z => n5097);
   U1932 : MUX21L port map( A => n26, B => n2501, S => n2416, Z => n5096);
   U1933 : MUX21L port map( A => n1096, B => n2501, S => n2417, Z => n5095);
   U1934 : MUX21L port map( A => n25, B => n2501, S => n2418, Z => n5094);
   U1935 : MUX21L port map( A => n2501, B => n1103, S => n2419, Z => n5093);
   U1936 : MUX21L port map( A => n2501, B => n32, S => n2420, Z => n5092);
   U1937 : MUX21L port map( A => n2501, B => n1102, S => n2421, Z => n5091);
   U1938 : MUX21L port map( A => n2501, B => n31, S => n2422, Z => n5090);
   U1939 : MUX21L port map( A => n1101, B => n2501, S => n2423, Z => n5089);
   U1940 : MUX21L port map( A => n30, B => n2501, S => n2424, Z => n5088);
   U1941 : MUX21L port map( A => n1100, B => n2501, S => n2425, Z => n5087);
   U1942 : MUX21L port map( A => n29, B => n2501, S => n2426, Z => n5086);
   U1943 : MUX21L port map( A => n2501, B => n1107, S => n2427, Z => n5085);
   U1944 : MUX21L port map( A => n2501, B => n36, S => n2428, Z => n5084);
   U1945 : MUX21L port map( A => n2501, B => n1106, S => n2429, Z => n5083);
   U1946 : MUX21L port map( A => n2501, B => n35, S => n2430, Z => n5082);
   U1947 : MUX21L port map( A => n1105, B => n2501, S => n2431, Z => n5081);
   U1948 : MUX21L port map( A => n34, B => n2501, S => n2432, Z => n5080);
   U1949 : MUX21L port map( A => n1104, B => n2501, S => n2433, Z => n5079);
   U1950 : MUX21L port map( A => n33, B => n2501, S => n2434, Z => n5078);
   U1951 : MUX21L port map( A => n2501, B => n1111, S => n2435, Z => n5077);
   U1952 : MUX21L port map( A => n2501, B => n40, S => n2436, Z => n5076);
   U1953 : MUX21L port map( A => n2501, B => n1110, S => n2437, Z => n5075);
   U1954 : MUX21L port map( A => n2501, B => n39, S => n2438, Z => n5074);
   U1955 : MUX21L port map( A => n1109, B => n2501, S => n2439, Z => n5073);
   U1956 : MUX21L port map( A => n38, B => n2501, S => n2440, Z => n5072);
   U1957 : MUX21L port map( A => n1108, B => n2501, S => n2441, Z => n5071);
   U1958 : MUX21L port map( A => n37, B => n2501, S => n2442, Z => n5070);
   U1959 : MUX21L port map( A => n2501, B => n1083, S => n2443, Z => n5069);
   U1960 : MUX21L port map( A => n2501, B => n12, S => n2444, Z => n5068);
   U1961 : MUX21L port map( A => n2501, B => n1082, S => n2445, Z => n5067);
   U1962 : MUX21L port map( A => n2501, B => n11, S => n2446, Z => n5066);
   U1963 : MUX21L port map( A => n1081, B => n2501, S => n2447, Z => n5065);
   U1964 : MUX21L port map( A => n10, B => n2501, S => n2448, Z => n5064);
   U1965 : MUX21L port map( A => n1080, B => n2501, S => n2449, Z => n5063);
   U1966 : MUX21L port map( A => n9, B => n2501, S => n2450, Z => n5062);
   U1967 : MUX21L port map( A => n2501, B => n1087, S => n2451, Z => n5061);
   U1968 : MUX21L port map( A => n2501, B => n16, S => n2452, Z => n5060);
   U1969 : MUX21L port map( A => n2501, B => n1086, S => n2453, Z => n5059);
   U1970 : MUX21L port map( A => n2501, B => n15, S => n2454, Z => n5058);
   U1971 : MUX21L port map( A => n1085, B => n2501, S => n2455, Z => n5057);
   U1972 : MUX21L port map( A => n14, B => n2501, S => n2456, Z => n5056);
   U1973 : MUX21L port map( A => n1084, B => n2501, S => n2457, Z => n5055);
   U1974 : MUX21L port map( A => n13, B => n2501, S => n2458, Z => n5054);
   U1975 : MUX21L port map( A => n2501, B => n1091, S => n2459, Z => n5053);
   U1976 : MUX21L port map( A => n2501, B => n20, S => n2460, Z => n5052);
   U1977 : MUX21L port map( A => n2501, B => n1090, S => n2461, Z => n5051);
   U1978 : MUX21L port map( A => n2501, B => n19, S => n2462, Z => n5050);
   U1979 : MUX21L port map( A => n1089, B => n2501, S => n2463, Z => n5049);
   U1980 : MUX21L port map( A => n18, B => n2501, S => n2464, Z => n5048);
   U1981 : MUX21L port map( A => n1088, B => n2501, S => n2465, Z => n5047);
   U1982 : MUX21L port map( A => n17, B => n2501, S => n2466, Z => n5046);
   U1983 : MUX21L port map( A => n2501, B => n1095, S => n2467, Z => n5045);
   U1984 : MUX21L port map( A => n2501, B => n24, S => n2468, Z => n5044);
   U1985 : MUX21L port map( A => n2501, B => n1094, S => n2469, Z => n5043);
   U1986 : MUX21L port map( A => n2501, B => n23, S => n2470, Z => n5042);
   U1987 : MUX21L port map( A => n1093, B => n2501, S => n2471, Z => n5041);
   U1988 : MUX21L port map( A => n22, B => n2501, S => n2472, Z => n5040);
   U1989 : MUX21L port map( A => n1092, B => n2501, S => n2473, Z => n5039);
   U1990 : MUX21L port map( A => n21, B => n2501, S => n2474, Z => n5038);
   U1991 : AO2 port map( A => v_TEMP_VECTOR_7_port, B => n2475, C => 
                           v_KEY32_IN_7_port, D => n2476, Z => n2501);
   U1992 : MUX21L port map( A => n2502, B => n1227, S => n2411, Z => n5037);
   U1993 : MUX21L port map( A => n2502, B => n156, S => n2412, Z => n5036);
   U1994 : MUX21L port map( A => n2502, B => n1226, S => n2413, Z => n5035);
   U1995 : MUX21L port map( A => n2502, B => n155, S => n2414, Z => n5034);
   U1996 : MUX21L port map( A => n1225, B => n2502, S => n2415, Z => n5033);
   U1997 : MUX21L port map( A => n154, B => n2502, S => n2416, Z => n5032);
   U1998 : MUX21L port map( A => n1224, B => n2502, S => n2417, Z => n5031);
   U1999 : MUX21L port map( A => n153, B => n2502, S => n2418, Z => n5030);
   U2000 : MUX21L port map( A => n2502, B => n1231, S => n2419, Z => n5029);
   U2001 : MUX21L port map( A => n2502, B => n160, S => n2420, Z => n5028);
   U2002 : MUX21L port map( A => n2502, B => n1230, S => n2421, Z => n5027);
   U2003 : MUX21L port map( A => n2502, B => n159, S => n2422, Z => n5026);
   U2004 : MUX21L port map( A => n1229, B => n2502, S => n2423, Z => n5025);
   U2005 : MUX21L port map( A => n158, B => n2502, S => n2424, Z => n5024);
   U2006 : MUX21L port map( A => n1228, B => n2502, S => n2425, Z => n5023);
   U2007 : MUX21L port map( A => n157, B => n2502, S => n2426, Z => n5022);
   U2008 : MUX21L port map( A => n2502, B => n1235, S => n2427, Z => n5021);
   U2009 : MUX21L port map( A => n2502, B => n164, S => n2428, Z => n5020);
   U2010 : MUX21L port map( A => n2502, B => n1234, S => n2429, Z => n5019);
   U2011 : MUX21L port map( A => n2502, B => n163, S => n2430, Z => n5018);
   U2012 : MUX21L port map( A => n1233, B => n2502, S => n2431, Z => n5017);
   U2013 : MUX21L port map( A => n162, B => n2502, S => n2432, Z => n5016);
   U2014 : MUX21L port map( A => n1232, B => n2502, S => n2433, Z => n5015);
   U2015 : MUX21L port map( A => n161, B => n2502, S => n2434, Z => n5014);
   U2016 : MUX21L port map( A => n2502, B => n1239, S => n2435, Z => n5013);
   U2017 : MUX21L port map( A => n2502, B => n168, S => n2436, Z => n5012);
   U2018 : MUX21L port map( A => n2502, B => n1238, S => n2437, Z => n5011);
   U2019 : MUX21L port map( A => n2502, B => n167, S => n2438, Z => n5010);
   U2020 : MUX21L port map( A => n1237, B => n2502, S => n2439, Z => n5009);
   U2021 : MUX21L port map( A => n166, B => n2502, S => n2440, Z => n5008);
   U2022 : MUX21L port map( A => n1236, B => n2502, S => n2441, Z => n5007);
   U2023 : MUX21L port map( A => n165, B => n2502, S => n2442, Z => n5006);
   U2024 : MUX21L port map( A => n2502, B => n1211, S => n2443, Z => n5005);
   U2025 : MUX21L port map( A => n2502, B => n140, S => n2444, Z => n5004);
   U2026 : MUX21L port map( A => n2502, B => n1210, S => n2445, Z => n5003);
   U2027 : MUX21L port map( A => n2502, B => n139, S => n2446, Z => n5002);
   U2028 : MUX21L port map( A => n1209, B => n2502, S => n2447, Z => n5001);
   U2029 : MUX21L port map( A => n138, B => n2502, S => n2448, Z => n5000);
   U2030 : MUX21L port map( A => n1208, B => n2502, S => n2449, Z => n4999);
   U2031 : MUX21L port map( A => n137, B => n2502, S => n2450, Z => n4998);
   U2032 : MUX21L port map( A => n2502, B => n1215, S => n2451, Z => n4997);
   U2033 : MUX21L port map( A => n2502, B => n144, S => n2452, Z => n4996);
   U2034 : MUX21L port map( A => n2502, B => n1214, S => n2453, Z => n4995);
   U2035 : MUX21L port map( A => n2502, B => n143, S => n2454, Z => n4994);
   U2036 : MUX21L port map( A => n1213, B => n2502, S => n2455, Z => n4993);
   U2037 : MUX21L port map( A => n142, B => n2502, S => n2456, Z => n4992);
   U2038 : MUX21L port map( A => n1212, B => n2502, S => n2457, Z => n4991);
   U2039 : MUX21L port map( A => n141, B => n2502, S => n2458, Z => n4990);
   U2040 : MUX21L port map( A => n2502, B => n1219, S => n2459, Z => n4989);
   U2041 : MUX21L port map( A => n2502, B => n148, S => n2460, Z => n4988);
   U2042 : MUX21L port map( A => n2502, B => n1218, S => n2461, Z => n4987);
   U2043 : MUX21L port map( A => n2502, B => n147, S => n2462, Z => n4986);
   U2044 : MUX21L port map( A => n1217, B => n2502, S => n2463, Z => n4985);
   U2045 : MUX21L port map( A => n146, B => n2502, S => n2464, Z => n4984);
   U2046 : MUX21L port map( A => n1216, B => n2502, S => n2465, Z => n4983);
   U2047 : MUX21L port map( A => n145, B => n2502, S => n2466, Z => n4982);
   U2048 : MUX21L port map( A => n2502, B => n1223, S => n2467, Z => n4981);
   U2049 : MUX21L port map( A => n2502, B => n152, S => n2468, Z => n4980);
   U2050 : MUX21L port map( A => n2502, B => n1222, S => n2469, Z => n4979);
   U2051 : MUX21L port map( A => n2502, B => n151, S => n2470, Z => n4978);
   U2052 : MUX21L port map( A => n1221, B => n2502, S => n2471, Z => n4977);
   U2053 : MUX21L port map( A => n150, B => n2502, S => n2472, Z => n4976);
   U2054 : MUX21L port map( A => n1220, B => n2502, S => n2473, Z => n4975);
   U2055 : MUX21L port map( A => n149, B => n2502, S => n2474, Z => n4974);
   U2056 : AO2 port map( A => v_TEMP_VECTOR_6_port, B => n2475, C => 
                           v_KEY32_IN_6_port, D => n2476, Z => n2502);
   U2057 : MUX21L port map( A => n2503, B => n1355, S => n2411, Z => n4973);
   U2058 : MUX21L port map( A => n2503, B => n284, S => n2412, Z => n4972);
   U2059 : MUX21L port map( A => n2503, B => n1354, S => n2413, Z => n4971);
   U2060 : MUX21L port map( A => n2503, B => n283, S => n2414, Z => n4970);
   U2061 : MUX21L port map( A => n1353, B => n2503, S => n2415, Z => n4969);
   U2062 : MUX21L port map( A => n282, B => n2503, S => n2416, Z => n4968);
   U2063 : MUX21L port map( A => n1352, B => n2503, S => n2417, Z => n4967);
   U2064 : MUX21L port map( A => n281, B => n2503, S => n2418, Z => n4966);
   U2065 : MUX21L port map( A => n2503, B => n1359, S => n2419, Z => n4965);
   U2066 : MUX21L port map( A => n2503, B => n288, S => n2420, Z => n4964);
   U2067 : MUX21L port map( A => n2503, B => n1358, S => n2421, Z => n4963);
   U2068 : MUX21L port map( A => n2503, B => n287, S => n2422, Z => n4962);
   U2069 : MUX21L port map( A => n1357, B => n2503, S => n2423, Z => n4961);
   U2070 : MUX21L port map( A => n286, B => n2503, S => n2424, Z => n4960);
   U2071 : MUX21L port map( A => n1356, B => n2503, S => n2425, Z => n4959);
   U2072 : MUX21L port map( A => n285, B => n2503, S => n2426, Z => n4958);
   U2073 : MUX21L port map( A => n2503, B => n1363, S => n2427, Z => n4957);
   U2074 : MUX21L port map( A => n2503, B => n292, S => n2428, Z => n4956);
   U2075 : MUX21L port map( A => n2503, B => n1362, S => n2429, Z => n4955);
   U2076 : MUX21L port map( A => n2503, B => n291, S => n2430, Z => n4954);
   U2077 : MUX21L port map( A => n1361, B => n2503, S => n2431, Z => n4953);
   U2078 : MUX21L port map( A => n290, B => n2503, S => n2432, Z => n4952);
   U2079 : MUX21L port map( A => n1360, B => n2503, S => n2433, Z => n4951);
   U2080 : MUX21L port map( A => n289, B => n2503, S => n2434, Z => n4950);
   U2081 : MUX21L port map( A => n2503, B => n1367, S => n2435, Z => n4949);
   U2082 : MUX21L port map( A => n2503, B => n296, S => n2436, Z => n4948);
   U2083 : MUX21L port map( A => n2503, B => n1366, S => n2437, Z => n4947);
   U2084 : MUX21L port map( A => n2503, B => n295, S => n2438, Z => n4946);
   U2085 : MUX21L port map( A => n1365, B => n2503, S => n2439, Z => n4945);
   U2086 : MUX21L port map( A => n294, B => n2503, S => n2440, Z => n4944);
   U2087 : MUX21L port map( A => n1364, B => n2503, S => n2441, Z => n4943);
   U2088 : MUX21L port map( A => n293, B => n2503, S => n2442, Z => n4942);
   U2089 : MUX21L port map( A => n2503, B => n1339, S => n2443, Z => n4941);
   U2090 : MUX21L port map( A => n2503, B => n268, S => n2444, Z => n4940);
   U2091 : MUX21L port map( A => n2503, B => n1338, S => n2445, Z => n4939);
   U2092 : MUX21L port map( A => n2503, B => n267, S => n2446, Z => n4938);
   U2093 : MUX21L port map( A => n1337, B => n2503, S => n2447, Z => n4937);
   U2094 : MUX21L port map( A => n266, B => n2503, S => n2448, Z => n4936);
   U2095 : MUX21L port map( A => n1336, B => n2503, S => n2449, Z => n4935);
   U2096 : MUX21L port map( A => n265, B => n2503, S => n2450, Z => n4934);
   U2097 : MUX21L port map( A => n2503, B => n1343, S => n2451, Z => n4933);
   U2098 : MUX21L port map( A => n2503, B => n272, S => n2452, Z => n4932);
   U2099 : MUX21L port map( A => n2503, B => n1342, S => n2453, Z => n4931);
   U2100 : MUX21L port map( A => n2503, B => n271, S => n2454, Z => n4930);
   U2101 : MUX21L port map( A => n1341, B => n2503, S => n2455, Z => n4929);
   U2102 : MUX21L port map( A => n270, B => n2503, S => n2456, Z => n4928);
   U2103 : MUX21L port map( A => n1340, B => n2503, S => n2457, Z => n4927);
   U2104 : MUX21L port map( A => n269, B => n2503, S => n2458, Z => n4926);
   U2105 : MUX21L port map( A => n2503, B => n1347, S => n2459, Z => n4925);
   U2106 : MUX21L port map( A => n2503, B => n276, S => n2460, Z => n4924);
   U2107 : MUX21L port map( A => n2503, B => n1346, S => n2461, Z => n4923);
   U2108 : MUX21L port map( A => n2503, B => n275, S => n2462, Z => n4922);
   U2109 : MUX21L port map( A => n1345, B => n2503, S => n2463, Z => n4921);
   U2110 : MUX21L port map( A => n274, B => n2503, S => n2464, Z => n4920);
   U2111 : MUX21L port map( A => n1344, B => n2503, S => n2465, Z => n4919);
   U2112 : MUX21L port map( A => n273, B => n2503, S => n2466, Z => n4918);
   U2113 : MUX21L port map( A => n2503, B => n1351, S => n2467, Z => n4917);
   U2114 : MUX21L port map( A => n2503, B => n280, S => n2468, Z => n4916);
   U2115 : MUX21L port map( A => n2503, B => n1350, S => n2469, Z => n4915);
   U2116 : MUX21L port map( A => n2503, B => n279, S => n2470, Z => n4914);
   U2117 : MUX21L port map( A => n1349, B => n2503, S => n2471, Z => n4913);
   U2118 : MUX21L port map( A => n278, B => n2503, S => n2472, Z => n4912);
   U2119 : MUX21L port map( A => n1348, B => n2503, S => n2473, Z => n4911);
   U2120 : MUX21L port map( A => n277, B => n2503, S => n2474, Z => n4910);
   U2121 : AO2 port map( A => v_TEMP_VECTOR_5_port, B => n2475, C => 
                           v_KEY32_IN_5_port, D => n2476, Z => n2503);
   U2122 : MUX21L port map( A => n2504, B => n1483, S => n2411, Z => n4909);
   U2123 : MUX21L port map( A => n2504, B => n412, S => n2412, Z => n4908);
   U2124 : MUX21L port map( A => n2504, B => n1482, S => n2413, Z => n4907);
   U2125 : MUX21L port map( A => n2504, B => n411, S => n2414, Z => n4906);
   U2126 : MUX21L port map( A => n1481, B => n2504, S => n2415, Z => n4905);
   U2127 : MUX21L port map( A => n410, B => n2504, S => n2416, Z => n4904);
   U2128 : MUX21L port map( A => n1480, B => n2504, S => n2417, Z => n4903);
   U2129 : MUX21L port map( A => n409, B => n2504, S => n2418, Z => n4902);
   U2130 : MUX21L port map( A => n2504, B => n1487, S => n2419, Z => n4901);
   U2131 : MUX21L port map( A => n2504, B => n416, S => n2420, Z => n4900);
   U2132 : MUX21L port map( A => n2504, B => n1486, S => n2421, Z => n4899);
   U2133 : MUX21L port map( A => n2504, B => n415, S => n2422, Z => n4898);
   U2134 : MUX21L port map( A => n1485, B => n2504, S => n2423, Z => n4897);
   U2135 : MUX21L port map( A => n414, B => n2504, S => n2424, Z => n4896);
   U2136 : MUX21L port map( A => n1484, B => n2504, S => n2425, Z => n4895);
   U2137 : MUX21L port map( A => n413, B => n2504, S => n2426, Z => n4894);
   U2138 : MUX21L port map( A => n2504, B => n1491, S => n2427, Z => n4893);
   U2139 : MUX21L port map( A => n2504, B => n420, S => n2428, Z => n4892);
   U2140 : MUX21L port map( A => n2504, B => n1490, S => n2429, Z => n4891);
   U2141 : MUX21L port map( A => n2504, B => n419, S => n2430, Z => n4890);
   U2142 : MUX21L port map( A => n1489, B => n2504, S => n2431, Z => n4889);
   U2143 : MUX21L port map( A => n418, B => n2504, S => n2432, Z => n4888);
   U2144 : MUX21L port map( A => n1488, B => n2504, S => n2433, Z => n4887);
   U2145 : MUX21L port map( A => n417, B => n2504, S => n2434, Z => n4886);
   U2146 : MUX21L port map( A => n2504, B => n1495, S => n2435, Z => n4885);
   U2147 : MUX21L port map( A => n2504, B => n424, S => n2436, Z => n4884);
   U2148 : MUX21L port map( A => n2504, B => n1494, S => n2437, Z => n4883);
   U2149 : MUX21L port map( A => n2504, B => n423, S => n2438, Z => n4882);
   U2150 : MUX21L port map( A => n1493, B => n2504, S => n2439, Z => n4881);
   U2151 : MUX21L port map( A => n422, B => n2504, S => n2440, Z => n4880);
   U2152 : MUX21L port map( A => n1492, B => n2504, S => n2441, Z => n4879);
   U2153 : MUX21L port map( A => n421, B => n2504, S => n2442, Z => n4878);
   U2154 : MUX21L port map( A => n2504, B => n1467, S => n2443, Z => n4877);
   U2155 : MUX21L port map( A => n2504, B => n396, S => n2444, Z => n4876);
   U2156 : MUX21L port map( A => n2504, B => n1466, S => n2445, Z => n4875);
   U2157 : MUX21L port map( A => n2504, B => n395, S => n2446, Z => n4874);
   U2158 : MUX21L port map( A => n1465, B => n2504, S => n2447, Z => n4873);
   U2159 : MUX21L port map( A => n394, B => n2504, S => n2448, Z => n4872);
   U2160 : MUX21L port map( A => n1464, B => n2504, S => n2449, Z => n4871);
   U2161 : MUX21L port map( A => n393, B => n2504, S => n2450, Z => n4870);
   U2162 : MUX21L port map( A => n2504, B => n1471, S => n2451, Z => n4869);
   U2163 : MUX21L port map( A => n2504, B => n400, S => n2452, Z => n4868);
   U2164 : MUX21L port map( A => n2504, B => n1470, S => n2453, Z => n4867);
   U2165 : MUX21L port map( A => n2504, B => n399, S => n2454, Z => n4866);
   U2166 : MUX21L port map( A => n1469, B => n2504, S => n2455, Z => n4865);
   U2167 : MUX21L port map( A => n398, B => n2504, S => n2456, Z => n4864);
   U2168 : MUX21L port map( A => n1468, B => n2504, S => n2457, Z => n4863);
   U2169 : MUX21L port map( A => n397, B => n2504, S => n2458, Z => n4862);
   U2170 : MUX21L port map( A => n2504, B => n1475, S => n2459, Z => n4861);
   U2171 : MUX21L port map( A => n2504, B => n404, S => n2460, Z => n4860);
   U2172 : MUX21L port map( A => n2504, B => n1474, S => n2461, Z => n4859);
   U2173 : MUX21L port map( A => n2504, B => n403, S => n2462, Z => n4858);
   U2174 : MUX21L port map( A => n1473, B => n2504, S => n2463, Z => n4857);
   U2175 : MUX21L port map( A => n402, B => n2504, S => n2464, Z => n4856);
   U2176 : MUX21L port map( A => n1472, B => n2504, S => n2465, Z => n4855);
   U2177 : MUX21L port map( A => n401, B => n2504, S => n2466, Z => n4854);
   U2178 : MUX21L port map( A => n2504, B => n1479, S => n2467, Z => n4853);
   U2179 : MUX21L port map( A => n2504, B => n408, S => n2468, Z => n4852);
   U2180 : MUX21L port map( A => n2504, B => n1478, S => n2469, Z => n4851);
   U2181 : MUX21L port map( A => n2504, B => n407, S => n2470, Z => n4850);
   U2182 : MUX21L port map( A => n1477, B => n2504, S => n2471, Z => n4849);
   U2183 : MUX21L port map( A => n406, B => n2504, S => n2472, Z => n4848);
   U2184 : MUX21L port map( A => n1476, B => n2504, S => n2473, Z => n4847);
   U2185 : MUX21L port map( A => n405, B => n2504, S => n2474, Z => n4846);
   U2186 : AO2 port map( A => v_TEMP_VECTOR_4_port, B => n2475, C => 
                           v_KEY32_IN_4_port, D => n2476, Z => n2504);
   U2187 : MUX21L port map( A => n2505, B => n1611, S => n2411, Z => n4845);
   U2188 : MUX21L port map( A => n2505, B => n540, S => n2412, Z => n4844);
   U2189 : MUX21L port map( A => n2505, B => n1610, S => n2413, Z => n4843);
   U2190 : MUX21L port map( A => n2505, B => n539, S => n2414, Z => n4842);
   U2191 : MUX21L port map( A => n1609, B => n2505, S => n2415, Z => n4841);
   U2192 : MUX21L port map( A => n538, B => n2505, S => n2416, Z => n4840);
   U2193 : MUX21L port map( A => n1608, B => n2505, S => n2417, Z => n4839);
   U2194 : MUX21L port map( A => n537, B => n2505, S => n2418, Z => n4838);
   U2195 : MUX21L port map( A => n2505, B => n1615, S => n2419, Z => n4837);
   U2196 : MUX21L port map( A => n2505, B => n544, S => n2420, Z => n4836);
   U2197 : MUX21L port map( A => n2505, B => n1614, S => n2421, Z => n4835);
   U2198 : MUX21L port map( A => n2505, B => n543, S => n2422, Z => n4834);
   U2199 : MUX21L port map( A => n1613, B => n2505, S => n2423, Z => n4833);
   U2200 : MUX21L port map( A => n542, B => n2505, S => n2424, Z => n4832);
   U2201 : MUX21L port map( A => n1612, B => n2505, S => n2425, Z => n4831);
   U2202 : MUX21L port map( A => n541, B => n2505, S => n2426, Z => n4830);
   U2203 : MUX21L port map( A => n2505, B => n1619, S => n2427, Z => n4829);
   U2204 : MUX21L port map( A => n2505, B => n548, S => n2428, Z => n4828);
   U2205 : MUX21L port map( A => n2505, B => n1618, S => n2429, Z => n4827);
   U2206 : MUX21L port map( A => n2505, B => n547, S => n2430, Z => n4826);
   U2207 : MUX21L port map( A => n1617, B => n2505, S => n2431, Z => n4825);
   U2208 : MUX21L port map( A => n546, B => n2505, S => n2432, Z => n4824);
   U2209 : MUX21L port map( A => n1616, B => n2505, S => n2433, Z => n4823);
   U2210 : MUX21L port map( A => n545, B => n2505, S => n2434, Z => n4822);
   U2211 : MUX21L port map( A => n2505, B => n1623, S => n2435, Z => n4821);
   U2212 : MUX21L port map( A => n2505, B => n552, S => n2436, Z => n4820);
   U2213 : MUX21L port map( A => n2505, B => n1622, S => n2437, Z => n4819);
   U2214 : MUX21L port map( A => n2505, B => n551, S => n2438, Z => n4818);
   U2215 : MUX21L port map( A => n1621, B => n2505, S => n2439, Z => n4817);
   U2216 : MUX21L port map( A => n550, B => n2505, S => n2440, Z => n4816);
   U2217 : MUX21L port map( A => n1620, B => n2505, S => n2441, Z => n4815);
   U2218 : MUX21L port map( A => n549, B => n2505, S => n2442, Z => n4814);
   U2219 : MUX21L port map( A => n2505, B => n1595, S => n2443, Z => n4813);
   U2220 : MUX21L port map( A => n2505, B => n524, S => n2444, Z => n4812);
   U2221 : MUX21L port map( A => n2505, B => n1594, S => n2445, Z => n4811);
   U2222 : MUX21L port map( A => n2505, B => n523, S => n2446, Z => n4810);
   U2223 : MUX21L port map( A => n1593, B => n2505, S => n2447, Z => n4809);
   U2224 : MUX21L port map( A => n522, B => n2505, S => n2448, Z => n4808);
   U2225 : MUX21L port map( A => n1592, B => n2505, S => n2449, Z => n4807);
   U2226 : MUX21L port map( A => n521, B => n2505, S => n2450, Z => n4806);
   U2227 : MUX21L port map( A => n2505, B => n1599, S => n2451, Z => n4805);
   U2228 : MUX21L port map( A => n2505, B => n528, S => n2452, Z => n4804);
   U2229 : MUX21L port map( A => n2505, B => n1598, S => n2453, Z => n4803);
   U2230 : MUX21L port map( A => n2505, B => n527, S => n2454, Z => n4802);
   U2231 : MUX21L port map( A => n1597, B => n2505, S => n2455, Z => n4801);
   U2232 : MUX21L port map( A => n526, B => n2505, S => n2456, Z => n4800);
   U2233 : MUX21L port map( A => n1596, B => n2505, S => n2457, Z => n4799);
   U2234 : MUX21L port map( A => n525, B => n2505, S => n2458, Z => n4798);
   U2235 : MUX21L port map( A => n2505, B => n1603, S => n2459, Z => n4797);
   U2236 : MUX21L port map( A => n2505, B => n532, S => n2460, Z => n4796);
   U2237 : MUX21L port map( A => n2505, B => n1602, S => n2461, Z => n4795);
   U2238 : MUX21L port map( A => n2505, B => n531, S => n2462, Z => n4794);
   U2239 : MUX21L port map( A => n1601, B => n2505, S => n2463, Z => n4793);
   U2240 : MUX21L port map( A => n530, B => n2505, S => n2464, Z => n4792);
   U2241 : MUX21L port map( A => n1600, B => n2505, S => n2465, Z => n4791);
   U2242 : MUX21L port map( A => n529, B => n2505, S => n2466, Z => n4790);
   U2243 : MUX21L port map( A => n2505, B => n1607, S => n2467, Z => n4789);
   U2244 : MUX21L port map( A => n2505, B => n536, S => n2468, Z => n4788);
   U2245 : MUX21L port map( A => n2505, B => n1606, S => n2469, Z => n4787);
   U2246 : MUX21L port map( A => n2505, B => n535, S => n2470, Z => n4786);
   U2247 : MUX21L port map( A => n1605, B => n2505, S => n2471, Z => n4785);
   U2248 : MUX21L port map( A => n534, B => n2505, S => n2472, Z => n4784);
   U2249 : MUX21L port map( A => n1604, B => n2505, S => n2473, Z => n4783);
   U2250 : MUX21L port map( A => n533, B => n2505, S => n2474, Z => n4782);
   U2251 : AO2 port map( A => v_TEMP_VECTOR_3_port, B => n2475, C => 
                           v_KEY32_IN_3_port, D => n2476, Z => n2505);
   U2252 : MUX21L port map( A => n2506, B => n1739, S => n2411, Z => n4781);
   U2253 : MUX21L port map( A => n2506, B => n668, S => n2412, Z => n4780);
   U2254 : MUX21L port map( A => n2506, B => n1738, S => n2413, Z => n4779);
   U2255 : MUX21L port map( A => n2506, B => n667, S => n2414, Z => n4778);
   U2256 : MUX21L port map( A => n1737, B => n2506, S => n2415, Z => n4777);
   U2257 : MUX21L port map( A => n666, B => n2506, S => n2416, Z => n4776);
   U2258 : MUX21L port map( A => n1736, B => n2506, S => n2417, Z => n4775);
   U2259 : MUX21L port map( A => n665, B => n2506, S => n2418, Z => n4774);
   U2260 : MUX21L port map( A => n2506, B => n1743, S => n2419, Z => n4773);
   U2261 : MUX21L port map( A => n2506, B => n672, S => n2420, Z => n4772);
   U2262 : MUX21L port map( A => n2506, B => n1742, S => n2421, Z => n4771);
   U2263 : MUX21L port map( A => n2506, B => n671, S => n2422, Z => n4770);
   U2264 : MUX21L port map( A => n1741, B => n2506, S => n2423, Z => n4769);
   U2265 : MUX21L port map( A => n670, B => n2506, S => n2424, Z => n4768);
   U2266 : MUX21L port map( A => n1740, B => n2506, S => n2425, Z => n4767);
   U2267 : MUX21L port map( A => n669, B => n2506, S => n2426, Z => n4766);
   U2268 : MUX21L port map( A => n2506, B => n1747, S => n2427, Z => n4765);
   U2269 : MUX21L port map( A => n2506, B => n676, S => n2428, Z => n4764);
   U2270 : MUX21L port map( A => n2506, B => n1746, S => n2429, Z => n4763);
   U2271 : MUX21L port map( A => n2506, B => n675, S => n2430, Z => n4762);
   U2272 : MUX21L port map( A => n1745, B => n2506, S => n2431, Z => n4761);
   U2273 : MUX21L port map( A => n674, B => n2506, S => n2432, Z => n4760);
   U2274 : MUX21L port map( A => n1744, B => n2506, S => n2433, Z => n4759);
   U2275 : MUX21L port map( A => n673, B => n2506, S => n2434, Z => n4758);
   U2276 : MUX21L port map( A => n2506, B => n1751, S => n2435, Z => n4757);
   U2277 : MUX21L port map( A => n2506, B => n680, S => n2436, Z => n4756);
   U2278 : MUX21L port map( A => n2506, B => n1750, S => n2437, Z => n4755);
   U2279 : MUX21L port map( A => n2506, B => n679, S => n2438, Z => n4754);
   U2280 : MUX21L port map( A => n1749, B => n2506, S => n2439, Z => n4753);
   U2281 : MUX21L port map( A => n678, B => n2506, S => n2440, Z => n4752);
   U2282 : MUX21L port map( A => n1748, B => n2506, S => n2441, Z => n4751);
   U2283 : MUX21L port map( A => n677, B => n2506, S => n2442, Z => n4750);
   U2284 : MUX21L port map( A => n2506, B => n1723, S => n2443, Z => n4749);
   U2285 : MUX21L port map( A => n2506, B => n652, S => n2444, Z => n4748);
   U2286 : MUX21L port map( A => n2506, B => n1722, S => n2445, Z => n4747);
   U2287 : MUX21L port map( A => n2506, B => n651, S => n2446, Z => n4746);
   U2288 : MUX21L port map( A => n1721, B => n2506, S => n2447, Z => n4745);
   U2289 : MUX21L port map( A => n650, B => n2506, S => n2448, Z => n4744);
   U2290 : MUX21L port map( A => n1720, B => n2506, S => n2449, Z => n4743);
   U2291 : MUX21L port map( A => n649, B => n2506, S => n2450, Z => n4742);
   U2292 : MUX21L port map( A => n2506, B => n1727, S => n2451, Z => n4741);
   U2293 : MUX21L port map( A => n2506, B => n656, S => n2452, Z => n4740);
   U2294 : MUX21L port map( A => n2506, B => n1726, S => n2453, Z => n4739);
   U2295 : MUX21L port map( A => n2506, B => n655, S => n2454, Z => n4738);
   U2296 : MUX21L port map( A => n1725, B => n2506, S => n2455, Z => n4737);
   U2297 : MUX21L port map( A => n654, B => n2506, S => n2456, Z => n4736);
   U2298 : MUX21L port map( A => n1724, B => n2506, S => n2457, Z => n4735);
   U2299 : MUX21L port map( A => n653, B => n2506, S => n2458, Z => n4734);
   U2300 : MUX21L port map( A => n2506, B => n1731, S => n2459, Z => n4733);
   U2301 : MUX21L port map( A => n2506, B => n660, S => n2460, Z => n4732);
   U2302 : MUX21L port map( A => n2506, B => n1730, S => n2461, Z => n4731);
   U2303 : MUX21L port map( A => n2506, B => n659, S => n2462, Z => n4730);
   U2304 : MUX21L port map( A => n1729, B => n2506, S => n2463, Z => n4729);
   U2305 : MUX21L port map( A => n658, B => n2506, S => n2464, Z => n4728);
   U2306 : MUX21L port map( A => n1728, B => n2506, S => n2465, Z => n4727);
   U2307 : MUX21L port map( A => n657, B => n2506, S => n2466, Z => n4726);
   U2308 : MUX21L port map( A => n2506, B => n1735, S => n2467, Z => n4725);
   U2309 : MUX21L port map( A => n2506, B => n664, S => n2468, Z => n4724);
   U2310 : MUX21L port map( A => n2506, B => n1734, S => n2469, Z => n4723);
   U2311 : MUX21L port map( A => n2506, B => n663, S => n2470, Z => n4722);
   U2312 : MUX21L port map( A => n1733, B => n2506, S => n2471, Z => n4721);
   U2313 : MUX21L port map( A => n662, B => n2506, S => n2472, Z => n4720);
   U2314 : MUX21L port map( A => n1732, B => n2506, S => n2473, Z => n4719);
   U2315 : MUX21L port map( A => n661, B => n2506, S => n2474, Z => n4718);
   U2316 : AO2 port map( A => v_TEMP_VECTOR_2_port, B => n2475, C => 
                           v_KEY32_IN_2_port, D => n2476, Z => n2506);
   U2317 : MUX21L port map( A => n2507, B => n1867, S => n2411, Z => n4717);
   U2318 : MUX21L port map( A => n2507, B => n796, S => n2412, Z => n4716);
   U2319 : MUX21L port map( A => n2507, B => n1866, S => n2413, Z => n4715);
   U2320 : MUX21L port map( A => n2507, B => n795, S => n2414, Z => n4714);
   U2321 : MUX21L port map( A => n1865, B => n2507, S => n2415, Z => n4713);
   U2322 : MUX21L port map( A => n794, B => n2507, S => n2416, Z => n4712);
   U2323 : MUX21L port map( A => n1864, B => n2507, S => n2417, Z => n4711);
   U2324 : MUX21L port map( A => n793, B => n2507, S => n2418, Z => n4710);
   U2325 : MUX21L port map( A => n2507, B => n1871, S => n2419, Z => n4709);
   U2326 : MUX21L port map( A => n2507, B => n800, S => n2420, Z => n4708);
   U2327 : MUX21L port map( A => n2507, B => n1870, S => n2421, Z => n4707);
   U2328 : MUX21L port map( A => n2507, B => n799, S => n2422, Z => n4706);
   U2329 : MUX21L port map( A => n1869, B => n2507, S => n2423, Z => n4705);
   U2330 : MUX21L port map( A => n798, B => n2507, S => n2424, Z => n4704);
   U2331 : MUX21L port map( A => n1868, B => n2507, S => n2425, Z => n4703);
   U2332 : MUX21L port map( A => n797, B => n2507, S => n2426, Z => n4702);
   U2333 : MUX21L port map( A => n2507, B => n1875, S => n2427, Z => n4701);
   U2334 : MUX21L port map( A => n2507, B => n804, S => n2428, Z => n4700);
   U2335 : MUX21L port map( A => n2507, B => n1874, S => n2429, Z => n4699);
   U2336 : MUX21L port map( A => n2507, B => n803, S => n2430, Z => n4698);
   U2337 : MUX21L port map( A => n1873, B => n2507, S => n2431, Z => n4697);
   U2338 : MUX21L port map( A => n802, B => n2507, S => n2432, Z => n4696);
   U2339 : MUX21L port map( A => n1872, B => n2507, S => n2433, Z => n4695);
   U2340 : MUX21L port map( A => n801, B => n2507, S => n2434, Z => n4694);
   U2341 : MUX21L port map( A => n2507, B => n1879, S => n2435, Z => n4693);
   U2342 : MUX21L port map( A => n2507, B => n808, S => n2436, Z => n4692);
   U2343 : MUX21L port map( A => n2507, B => n1878, S => n2437, Z => n4691);
   U2344 : MUX21L port map( A => n2507, B => n807, S => n2438, Z => n4690);
   U2345 : MUX21L port map( A => n1877, B => n2507, S => n2439, Z => n4689);
   U2346 : MUX21L port map( A => n806, B => n2507, S => n2440, Z => n4688);
   U2347 : MUX21L port map( A => n1876, B => n2507, S => n2441, Z => n4687);
   U2348 : MUX21L port map( A => n805, B => n2507, S => n2442, Z => n4686);
   U2349 : MUX21L port map( A => n2507, B => n1851, S => n2443, Z => n4685);
   U2350 : MUX21L port map( A => n2507, B => n780, S => n2444, Z => n4684);
   U2351 : MUX21L port map( A => n2507, B => n1850, S => n2445, Z => n4683);
   U2352 : MUX21L port map( A => n2507, B => n779, S => n2446, Z => n4682);
   U2353 : MUX21L port map( A => n1849, B => n2507, S => n2447, Z => n4681);
   U2354 : MUX21L port map( A => n778, B => n2507, S => n2448, Z => n4680);
   U2355 : MUX21L port map( A => n1848, B => n2507, S => n2449, Z => n4679);
   U2356 : MUX21L port map( A => n777, B => n2507, S => n2450, Z => n4678);
   U2357 : MUX21L port map( A => n2507, B => n1855, S => n2451, Z => n4677);
   U2358 : MUX21L port map( A => n2507, B => n784, S => n2452, Z => n4676);
   U2359 : MUX21L port map( A => n2507, B => n1854, S => n2453, Z => n4675);
   U2360 : MUX21L port map( A => n2507, B => n783, S => n2454, Z => n4674);
   U2361 : MUX21L port map( A => n1853, B => n2507, S => n2455, Z => n4673);
   U2362 : MUX21L port map( A => n782, B => n2507, S => n2456, Z => n4672);
   U2363 : MUX21L port map( A => n1852, B => n2507, S => n2457, Z => n4671);
   U2364 : MUX21L port map( A => n781, B => n2507, S => n2458, Z => n4670);
   U2365 : MUX21L port map( A => n2507, B => n1859, S => n2459, Z => n4669);
   U2366 : MUX21L port map( A => n2507, B => n788, S => n2460, Z => n4668);
   U2367 : MUX21L port map( A => n2507, B => n1858, S => n2461, Z => n4667);
   U2368 : MUX21L port map( A => n2507, B => n787, S => n2462, Z => n4666);
   U2369 : MUX21L port map( A => n1857, B => n2507, S => n2463, Z => n4665);
   U2370 : MUX21L port map( A => n786, B => n2507, S => n2464, Z => n4664);
   U2371 : MUX21L port map( A => n1856, B => n2507, S => n2465, Z => n4663);
   U2372 : MUX21L port map( A => n785, B => n2507, S => n2466, Z => n4662);
   U2373 : MUX21L port map( A => n2507, B => n1863, S => n2467, Z => n4661);
   U2374 : MUX21L port map( A => n2507, B => n792, S => n2468, Z => n4660);
   U2375 : MUX21L port map( A => n2507, B => n1862, S => n2469, Z => n4659);
   U2376 : MUX21L port map( A => n2507, B => n791, S => n2470, Z => n4658);
   U2377 : MUX21L port map( A => n1861, B => n2507, S => n2471, Z => n4657);
   U2378 : MUX21L port map( A => n790, B => n2507, S => n2472, Z => n4656);
   U2379 : MUX21L port map( A => n1860, B => n2507, S => n2473, Z => n4655);
   U2380 : MUX21L port map( A => n789, B => n2507, S => n2474, Z => n4654);
   U2381 : AO2 port map( A => v_TEMP_VECTOR_1_port, B => n2475, C => 
                           v_KEY32_IN_1_port, D => n2476, Z => n2507);
   U2382 : MUX21L port map( A => n2508, B => n1995, S => n2411, Z => n4653);
   U2383 : ND2 port map( A => n2509, B => n2206, Z => n2411);
   U2384 : MUX21L port map( A => n2508, B => n924, S => n2412, Z => n4652);
   U2385 : ND2 port map( A => n2510, B => n2509, Z => n2412);
   U2386 : MUX21L port map( A => n2508, B => n1994, S => n2413, Z => n4651);
   U2387 : ND2 port map( A => n2511, B => n2509, Z => n2413);
   U2388 : MUX21L port map( A => n2508, B => n923, S => n2414, Z => n4650);
   U2389 : ND2 port map( A => n2512, B => n2509, Z => n2414);
   U2390 : IV port map( A => n2513, Z => n2509);
   U2391 : MUX21L port map( A => n1993, B => n2508, S => n2415, Z => n4649);
   U2392 : NR2 port map( A => n2513, B => n2202, Z => n2415);
   U2393 : MUX21L port map( A => n922, B => n2508, S => n2416, Z => n4648);
   U2394 : NR2 port map( A => n2514, B => n2513, Z => n2416);
   U2395 : MUX21L port map( A => n1992, B => n2508, S => n2417, Z => n4647);
   U2396 : NR2 port map( A => n2515, B => n2513, Z => n2417);
   U2397 : MUX21L port map( A => n921, B => n2508, S => n2418, Z => n4646);
   U2398 : NR2 port map( A => n2516, B => n2513, Z => n2418);
   U2399 : ND3 port map( A => n2, B => n1035, C => n2517, Z => n2513);
   U2400 : MUX21L port map( A => n2508, B => n1999, S => n2419, Z => n4645);
   U2401 : ND2 port map( A => n2518, B => n2206, Z => n2419);
   U2402 : MUX21L port map( A => n2508, B => n928, S => n2420, Z => n4644);
   U2403 : ND2 port map( A => n2518, B => n2510, Z => n2420);
   U2404 : MUX21L port map( A => n2508, B => n1998, S => n2421, Z => n4643);
   U2405 : ND2 port map( A => n2518, B => n2511, Z => n2421);
   U2406 : MUX21L port map( A => n2508, B => n927, S => n2422, Z => n4642);
   U2407 : ND2 port map( A => n2518, B => n2512, Z => n2422);
   U2408 : IV port map( A => n2519, Z => n2518);
   U2409 : MUX21L port map( A => n1997, B => n2508, S => n2423, Z => n4641);
   U2410 : NR2 port map( A => n2519, B => n2202, Z => n2423);
   U2411 : MUX21L port map( A => n926, B => n2508, S => n2424, Z => n4640);
   U2412 : NR2 port map( A => n2519, B => n2514, Z => n2424);
   U2413 : MUX21L port map( A => n1996, B => n2508, S => n2425, Z => n4639);
   U2414 : NR2 port map( A => n2519, B => n2515, Z => n2425);
   U2415 : MUX21L port map( A => n925, B => n2508, S => n2426, Z => n4638);
   U2416 : NR2 port map( A => n2519, B => n2516, Z => n2426);
   U2417 : ND3 port map( A => n6640, B => n2, C => n2517, Z => n2519);
   U2418 : MUX21L port map( A => n2508, B => n2003, S => n2427, Z => n4637);
   U2419 : ND2 port map( A => n2520, B => n2206, Z => n2427);
   U2420 : MUX21L port map( A => n2508, B => n932, S => n2428, Z => n4636);
   U2421 : ND2 port map( A => n2520, B => n2510, Z => n2428);
   U2422 : MUX21L port map( A => n2508, B => n2002, S => n2429, Z => n4635);
   U2423 : ND2 port map( A => n2520, B => n2511, Z => n2429);
   U2424 : MUX21L port map( A => n2508, B => n931, S => n2430, Z => n4634);
   U2425 : ND2 port map( A => n2520, B => n2512, Z => n2430);
   U2426 : IV port map( A => n2521, Z => n2520);
   U2427 : MUX21L port map( A => n2001, B => n2508, S => n2431, Z => n4633);
   U2428 : NR2 port map( A => n2521, B => n2202, Z => n2431);
   U2429 : MUX21L port map( A => n930, B => n2508, S => n2432, Z => n4632);
   U2430 : NR2 port map( A => n2521, B => n2514, Z => n2432);
   U2431 : MUX21L port map( A => n2000, B => n2508, S => n2433, Z => n4631);
   U2432 : NR2 port map( A => n2521, B => n2515, Z => n2433);
   U2433 : MUX21L port map( A => n929, B => n2508, S => n2434, Z => n4630);
   U2434 : NR2 port map( A => n2521, B => n2516, Z => n2434);
   U2435 : ND3 port map( A => n6639, B => n1035, C => n2517, Z => n2521);
   U2436 : MUX21L port map( A => n2508, B => n2007, S => n2435, Z => n4629);
   U2437 : ND2 port map( A => n2522, B => n2206, Z => n2435);
   U2438 : MUX21L port map( A => n2508, B => n936, S => n2436, Z => n4628);
   U2439 : ND2 port map( A => n2522, B => n2510, Z => n2436);
   U2440 : MUX21L port map( A => n2508, B => n2006, S => n2437, Z => n4627);
   U2441 : ND2 port map( A => n2522, B => n2511, Z => n2437);
   U2442 : MUX21L port map( A => n2508, B => n935, S => n2438, Z => n4626);
   U2443 : ND2 port map( A => n2522, B => n2512, Z => n2438);
   U2444 : IV port map( A => n2523, Z => n2522);
   U2445 : MUX21L port map( A => n2005, B => n2508, S => n2439, Z => n4625);
   U2446 : NR2 port map( A => n2523, B => n2202, Z => n2439);
   U2447 : MUX21L port map( A => n934, B => n2508, S => n2440, Z => n4624);
   U2448 : NR2 port map( A => n2523, B => n2514, Z => n2440);
   U2449 : MUX21L port map( A => n2004, B => n2508, S => n2441, Z => n4623);
   U2450 : NR2 port map( A => n2523, B => n2515, Z => n2441);
   U2451 : MUX21L port map( A => n933, B => n2508, S => n2442, Z => n4622);
   U2452 : NR2 port map( A => n2523, B => n2516, Z => n2442);
   U2453 : ND3 port map( A => n6639, B => n6640, C => n2517, Z => n2523);
   U2454 : NR3 port map( A => n2140, B => n6638, C => n1076, Z => n2517);
   U2455 : MUX21L port map( A => n2508, B => n1979, S => n2443, Z => n4621);
   U2456 : ND2 port map( A => n2524, B => n2206, Z => n2443);
   U2457 : MUX21L port map( A => n2508, B => n908, S => n2444, Z => n4620);
   U2458 : ND2 port map( A => n2524, B => n2510, Z => n2444);
   U2459 : MUX21L port map( A => n2508, B => n1978, S => n2445, Z => n4619);
   U2460 : ND2 port map( A => n2524, B => n2511, Z => n2445);
   U2461 : MUX21L port map( A => n2508, B => n907, S => n2446, Z => n4618);
   U2462 : ND2 port map( A => n2524, B => n2512, Z => n2446);
   U2463 : IV port map( A => n2525, Z => n2524);
   U2464 : MUX21L port map( A => n1977, B => n2508, S => n2447, Z => n4617);
   U2465 : NR2 port map( A => n2525, B => n2202, Z => n2447);
   U2466 : MUX21L port map( A => n906, B => n2508, S => n2448, Z => n4616);
   U2467 : NR2 port map( A => n2525, B => n2514, Z => n2448);
   U2468 : MUX21L port map( A => n1976, B => n2508, S => n2449, Z => n4615);
   U2469 : NR2 port map( A => n2525, B => n2515, Z => n2449);
   U2470 : MUX21L port map( A => n905, B => n2508, S => n2450, Z => n4614);
   U2471 : NR2 port map( A => n2525, B => n2516, Z => n2450);
   U2472 : ND3 port map( A => n2, B => n1035, C => n2526, Z => n2525);
   U2473 : MUX21L port map( A => n2508, B => n1983, S => n2451, Z => n4613);
   U2474 : ND2 port map( A => n2527, B => n2206, Z => n2451);
   U2475 : MUX21L port map( A => n2508, B => n912, S => n2452, Z => n4612);
   U2476 : ND2 port map( A => n2527, B => n2510, Z => n2452);
   U2477 : MUX21L port map( A => n2508, B => n1982, S => n2453, Z => n4611);
   U2478 : ND2 port map( A => n2527, B => n2511, Z => n2453);
   U2479 : MUX21L port map( A => n2508, B => n911, S => n2454, Z => n4610);
   U2480 : ND2 port map( A => n2527, B => n2512, Z => n2454);
   U2481 : IV port map( A => n2528, Z => n2527);
   U2482 : MUX21L port map( A => n1981, B => n2508, S => n2455, Z => n4609);
   U2483 : NR2 port map( A => n2528, B => n2202, Z => n2455);
   U2484 : MUX21L port map( A => n910, B => n2508, S => n2456, Z => n4608);
   U2485 : NR2 port map( A => n2528, B => n2514, Z => n2456);
   U2486 : MUX21L port map( A => n1980, B => n2508, S => n2457, Z => n4607);
   U2487 : NR2 port map( A => n2528, B => n2515, Z => n2457);
   U2488 : MUX21L port map( A => n909, B => n2508, S => n2458, Z => n4606);
   U2489 : NR2 port map( A => n2528, B => n2516, Z => n2458);
   U2490 : ND3 port map( A => n6640, B => n2, C => n2526, Z => n2528);
   U2491 : MUX21L port map( A => n2508, B => n1987, S => n2459, Z => n4605);
   U2492 : ND2 port map( A => n2529, B => n2206, Z => n2459);
   U2493 : MUX21L port map( A => n2508, B => n916, S => n2460, Z => n4604);
   U2494 : ND2 port map( A => n2529, B => n2510, Z => n2460);
   U2495 : MUX21L port map( A => n2508, B => n1986, S => n2461, Z => n4603);
   U2496 : ND2 port map( A => n2529, B => n2511, Z => n2461);
   U2497 : MUX21L port map( A => n2508, B => n915, S => n2462, Z => n4602);
   U2498 : ND2 port map( A => n2529, B => n2512, Z => n2462);
   U2499 : IV port map( A => n2530, Z => n2529);
   U2500 : MUX21L port map( A => n1985, B => n2508, S => n2463, Z => n4601);
   U2501 : NR2 port map( A => n2530, B => n2202, Z => n2463);
   U2502 : MUX21L port map( A => n914, B => n2508, S => n2464, Z => n4600);
   U2503 : NR2 port map( A => n2530, B => n2514, Z => n2464);
   U2504 : MUX21L port map( A => n1984, B => n2508, S => n2465, Z => n4599);
   U2505 : NR2 port map( A => n2530, B => n2515, Z => n2465);
   U2506 : MUX21L port map( A => n913, B => n2508, S => n2466, Z => n4598);
   U2507 : NR2 port map( A => n2530, B => n2516, Z => n2466);
   U2508 : ND3 port map( A => n6639, B => n1035, C => n2526, Z => n2530);
   U2509 : MUX21L port map( A => n2508, B => n1991, S => n2467, Z => n4597);
   U2510 : ND2 port map( A => n2531, B => n2206, Z => n2467);
   U2511 : NR3 port map( A => n6643, B => n6642, C => n6641, Z => n2206);
   U2512 : MUX21L port map( A => n2508, B => n920, S => n2468, Z => n4596);
   U2513 : ND2 port map( A => n2531, B => n2510, Z => n2468);
   U2514 : NR3 port map( A => n6641, B => n6642, C => n4, Z => n2510);
   U2515 : MUX21L port map( A => n2508, B => n1990, S => n2469, Z => n4595);
   U2516 : ND2 port map( A => n2531, B => n2511, Z => n2469);
   U2517 : NR2 port map( A => n2200, B => n6641, Z => n2511);
   U2518 : MUX21L port map( A => n2508, B => n919, S => n2470, Z => n4594);
   U2519 : ND2 port map( A => n2531, B => n2512, Z => n2470);
   U2520 : NR3 port map( A => n4, B => n6641, C => n1038, Z => n2512);
   U2521 : IV port map( A => n2532, Z => n2531);
   U2522 : MUX21L port map( A => n1989, B => n2508, S => n2471, Z => n4593);
   U2523 : NR2 port map( A => n2532, B => n2202, Z => n2471);
   U2524 : ND3 port map( A => n1038, B => n4, C => n6641, Z => n2202);
   U2525 : MUX21L port map( A => n918, B => n2508, S => n2472, Z => n4592);
   U2526 : NR2 port map( A => n2532, B => n2514, Z => n2472);
   U2527 : ND3 port map( A => n6643, B => n1038, C => n6641, Z => n2514);
   U2528 : MUX21L port map( A => n1988, B => n2508, S => n2473, Z => n4591);
   U2529 : NR2 port map( A => n2532, B => n2515, Z => n2473);
   U2530 : ND2 port map( A => n6641, B => n2533, Z => n2515);
   U2531 : IV port map( A => n2200, Z => n2533);
   U2532 : ND2 port map( A => n6642, B => n4, Z => n2200);
   U2533 : MUX21L port map( A => n917, B => n2508, S => n2474, Z => n4590);
   U2534 : NR2 port map( A => n2532, B => n2516, Z => n2474);
   U2535 : ND3 port map( A => n6642, B => n6643, C => n6641, Z => n2516);
   U2536 : ND3 port map( A => n6639, B => n6640, C => n2526, Z => n2532);
   U2537 : AN3 port map( A => n4470, B => CE_I, C => n6638, Z => n2526);
   U2538 : AO2 port map( A => v_TEMP_VECTOR_0_port, B => n2475, C => 
                           v_KEY32_IN_0_port, D => n2476, Z => n2508);
   U2539 : NR2 port map( A => n2534, B => n2476, Z => n2475);
   U2540 : AN3 port map( A => n1039, B => n6, C => n4469, Z => n2476);
   U2541 : IV port map( A => n2535, Z => n2534);
   U2542 : AO3 port map( A => n2390, B => n2189, C => n2536, D => n2409, Z => 
                           n2535);
   U2543 : ND2 port map( A => n2537, B => n2396, Z => n2409);
   U2544 : ND2 port map( A => n2396, B => n2538, Z => n2536);
   U2545 : AO7 port map( A => v_CALCULATION_CNTR_2_port, B => n7, C => n2539, Z
                           => n2538);
   U2546 : NR3 port map( A => n2540, B => v_CALCULATION_CNTR_3_port, C => n8, Z
                           => n2396);
   U2547 : AO6 port map( A => n1036, B => n2395, C => n2541, Z => n2390);
   U2548 : AO7 port map( A => CE_I, B => n1040, C => n2138, Z => n4589);
   U2549 : ND2 port map( A => VALID_KEY_I, B => CE_I, Z => n2138);
   U2550 : AO3 port map( A => n2542, B => n2543, C => n2544, D => n2545, Z => 
                           n4588);
   U2551 : AO2 port map( A => n2546, B => n2547, C => v_SUB_WORD_7_port, D => 
                           n2140, Z => n2545);
   U2552 : AO3 port map( A => n2548, B => n2549, C => n2550, D => n2551, Z => 
                           n2547);
   U2553 : AO1 port map( A => n2552, B => n2553, C => n2554, D => n2555, Z => 
                           n2551);
   U2554 : IV port map( A => n2556, Z => n2555);
   U2555 : AO4 port map( A => n2557, B => n2558, C => n2559, D => n2560, Z => 
                           n2554);
   U2556 : AO6 port map( A => n2561, B => n2562, C => n2563, Z => n2559);
   U2557 : NR2 port map( A => n2564, B => n2565, Z => n2557);
   U2558 : NR2 port map( A => n2566, B => n2567, Z => n2552);
   U2559 : AO2 port map( A => n2568, B => n2569, C => n2570, D => n2571, Z => 
                           n2550);
   U2560 : ND2 port map( A => n2572, B => n2573, Z => n2569);
   U2561 : IV port map( A => n2574, Z => n2548);
   U2562 : ND3 port map( A => n2575, B => n2576, C => n2577, Z => n2544);
   U2563 : MUX21L port map( A => n2578, B => n2579, S => n2580, Z => n2577);
   U2564 : AO1 port map( A => n2581, B => n2582, C => n2583, D => n2584, Z => 
                           n2579);
   U2565 : AO3 port map( A => n2585, B => n2586, C => n2587, D => n2588, Z => 
                           n2583);
   U2566 : OR3 port map( A => n2589, B => n2590, C => n2591, Z => n2588);
   U2567 : ND3 port map( A => n2592, B => n2593, C => n2594, Z => n2587);
   U2568 : AO3 port map( A => n2595, B => n2596, C => n2597, D => n2598, Z => 
                           n2578);
   U2569 : AO6 port map( A => n2599, B => n2600, C => n2601, Z => n2598);
   U2570 : AO4 port map( A => n2602, B => n2603, C => n2604, D => n2605, Z => 
                           n2601);
   U2571 : EO1 port map( A => n2606, B => n2584, C => n2607, D => n2558, Z => 
                           n2597);
   U2572 : AO3 port map( A => n2608, B => n2591, C => n2609, D => n2610, Z => 
                           n2606);
   U2573 : AO2 port map( A => n2611, B => n2612, C => n2613, D => n2614, Z => 
                           n2610);
   U2574 : AO7 port map( A => n2615, B => n2616, C => n2594, Z => n2609);
   U2575 : AN2 port map( A => n2573, B => n2617, Z => n2608);
   U2576 : AO3 port map( A => n2618, B => n2591, C => n2619, D => n2620, Z => 
                           n2576);
   U2577 : AO6 port map( A => n2594, B => n2621, C => n2622, Z => n2620);
   U2578 : EON1 port map( A => n2595, B => n2585, C => n2623, D => n2612, Z => 
                           n2622);
   U2579 : AN2 port map( A => n2624, B => n2625, Z => n2618);
   U2580 : AO3 port map( A => n2626, B => n2627, C => n2628, D => n2629, Z => 
                           n2543);
   U2581 : ND2 port map( A => n2630, B => n2553, Z => n2628);
   U2582 : AO3 port map( A => n2631, B => n2632, C => n2633, D => n2634, Z => 
                           n2542);
   U2583 : AO3 port map( A => n2591, B => n2635, C => n2636, D => n2637, Z => 
                           n2634);
   U2584 : AO1 port map( A => n2612, B => n2572, C => n2638, D => n2639, Z => 
                           n2637);
   U2585 : AO6 port map( A => n2640, B => n2641, C => n2642, Z => n2639);
   U2586 : NR2 port map( A => n2643, B => n2585, Z => n2638);
   U2587 : OR3 port map( A => n2566, B => n2644, C => n2645, Z => n2633);
   U2588 : IV port map( A => n2646, Z => n2631);
   U2589 : AO3 port map( A => CE_I, B => n1041, C => n2647, D => n2648, Z => 
                           n4587);
   U2590 : AO2 port map( A => n2649, B => n2650, C => n2651, D => n2652, Z => 
                           n2648);
   U2591 : AO1 port map( A => n2653, B => n2654, C => n2655, D => n2656, Z => 
                           n2652);
   U2592 : AO4 port map( A => n2657, B => n2658, C => n2659, D => n2626, Z => 
                           n2656);
   U2593 : AN2 port map( A => n2660, B => n2661, Z => n2659);
   U2594 : NR2 port map( A => n2662, B => n2611, Z => n2657);
   U2595 : EON1 port map( A => n2558, B => n2646, C => n2663, D => n2563, Z => 
                           n2655);
   U2596 : AO1 port map( A => n2599, B => n2664, C => n2665, D => n2666, Z => 
                           n2651);
   U2597 : AO4 port map( A => n2632, B => n2667, C => n2668, D => n2669, Z => 
                           n2665);
   U2598 : AO1 port map( A => n2670, B => n2553, C => n2671, D => n2672, Z => 
                           n2650);
   U2599 : NR2 port map( A => n2585, B => n2573, Z => n2672);
   U2600 : AO4 port map( A => n2621, B => n2596, C => n2626, D => n2663, Z => 
                           n2671);
   U2601 : NR4 port map( A => n2673, B => n2674, C => n2675, D => n2676, Z => 
                           n2649);
   U2602 : MUX21L port map( A => n2645, B => n2668, S => n2677, Z => n2676);
   U2603 : NR2 port map( A => n2632, B => n2678, Z => n2673);
   U2604 : OR3 port map( A => n2679, B => n2680, C => n2681, Z => n2647);
   U2605 : MUX21L port map( A => n2682, B => n2683, S => n2580, Z => n2681);
   U2606 : AO3 port map( A => n2684, B => n2642, C => n2636, D => n2685, Z => 
                           n2683);
   U2607 : AO1 port map( A => n2612, B => n2627, C => n2686, D => n2687, Z => 
                           n2685);
   U2608 : AN3 port map( A => n2688, B => n2593, C => n2595, Z => n2687);
   U2609 : AN3 port map( A => n2667, B => n2572, C => n2614, Z => n2686);
   U2610 : NR3 port map( A => n2689, B => n2690, C => n2691, Z => n2682);
   U2611 : AO4 port map( A => n2658, B => n2625, C => n2692, D => n2693, Z => 
                           n2691);
   U2612 : AO4 port map( A => n2626, B => n2694, C => n2643, D => n2645, Z => 
                           n2690);
   U2613 : AO3 port map( A => n2695, B => n2558, C => n2696, D => n2697, Z => 
                           n2689);
   U2614 : AO2 port map( A => n2698, B => n2699, C => n2700, D => n2599, Z => 
                           n2697);
   U2615 : ND2 port map( A => n2624, B => n2572, Z => n2699);
   U2616 : NR2 port map( A => n2566, B => n2701, Z => n2695);
   U2617 : AO1 port map( A => n2702, B => n2594, C => n2703, D => n2704, Z => 
                           n2679);
   U2618 : AO3 port map( A => n2705, B => n2585, C => n2706, D => n2707, Z => 
                           n2703);
   U2619 : ND3 port map( A => n2592, B => n2593, C => n2688, Z => n2707);
   U2620 : AO7 port map( A => n2611, B => n2590, C => n2612, Z => n2706);
   U2621 : AO3 port map( A => n2708, B => n2666, C => n2709, D => n2710, Z => 
                           n4586);
   U2622 : AO2 port map( A => n2711, B => n2712, C => n2140, D => n2105, Z => 
                           n2710);
   U2623 : AO3 port map( A => n2713, B => n2658, C => n2714, D => n2715, Z => 
                           n2712);
   U2624 : AO1 port map( A => n2716, B => n2717, C => n2718, D => n2719, Z => 
                           n2715);
   U2625 : AO6 port map( A => n2645, B => n2720, C => n2581, Z => n2719);
   U2626 : AO7 port map( A => n2677, B => n2721, C => n2561, Z => n2720);
   U2627 : IV port map( A => n2722, Z => n2677);
   U2628 : EON1 port map( A => n2723, B => n2603, C => n2568, D => n2724, Z => 
                           n2718);
   U2629 : AO2 port map( A => n2599, B => n2611, C => n2725, D => n2726, Z => 
                           n2714);
   U2630 : AO2 port map( A => n2727, B => n2728, C => n2729, D => n2730, Z => 
                           n2709);
   U2631 : ND4 port map( A => n2731, B => n2732, C => n2733, D => n2734, Z => 
                           n2730);
   U2632 : AO2 port map( A => n2735, B => n2698, C => n2563, D => n2560, Z => 
                           n2734);
   U2633 : NR2 port map( A => n2565, B => n2736, Z => n2735);
   U2634 : AO2 port map( A => n2570, B => n2627, C => n2725, D => n2641, Z => 
                           n2733);
   U2635 : MUX21L port map( A => n2737, B => n2738, S => n2739, Z => n2732);
   U2636 : NR2 port map( A => n2740, B => n2741, Z => n2738);
   U2637 : NR2 port map( A => n2664, B => n2658, Z => n2737);
   U2638 : AO2 port map( A => n2568, B => n2595, C => n2564, D => n2599, Z => 
                           n2731);
   U2639 : AO1 port map( A => n2698, B => n2616, C => n2742, D => n2743, Z => 
                           n2728);
   U2640 : NR3 port map( A => n2658, B => n2744, C => n2566, Z => n2743);
   U2641 : AN3 port map( A => n2636, B => n2745, C => n2746, Z => n2742);
   U2642 : AO2 port map( A => n2747, B => n2635, C => n2614, D => n2713, Z => 
                           n2746);
   U2643 : AO7 port map( A => n2748, B => n2694, C => n2692, Z => n2747);
   U2644 : AO1 port map( A => n2716, B => n2600, C => n2674, D => n2749, Z => 
                           n2727);
   U2645 : AO6 port map( A => n2625, B => n2592, C => n2645, Z => n2749);
   U2646 : AO1 port map( A => n2750, B => n2563, C => n2751, D => n2752, Z => 
                           n2708);
   U2647 : AO4 port map( A => n2670, B => n2668, C => n2558, D => n2753, Z => 
                           n2752);
   U2648 : IV port map( A => n2754, Z => n2670);
   U2649 : AO3 port map( A => n2755, B => n2658, C => n2756, D => n2757, Z => 
                           n2751);
   U2650 : AO2 port map( A => n2758, B => n2624, C => n2599, D => n2759, Z => 
                           n2757);
   U2651 : ND2 port map( A => n2722, B => n2760, Z => n2759);
   U2652 : AO7 port map( A => n2761, B => n2632, C => n2603, Z => n2758);
   U2653 : IV port map( A => n2762, Z => n2761);
   U2654 : OR3 port map( A => n2595, B => n2736, C => n2626, Z => n2756);
   U2655 : AN2 port map( A => n2660, B => n2669, Z => n2755);
   U2656 : ND3 port map( A => n2763, B => n2764, C => n2765, Z => n4585);
   U2657 : AO2 port map( A => n2766, B => n2767, C => n2140, D => n2106, Z => 
                           n2765);
   U2658 : AO1 port map( A => n2698, B => n2572, C => n2768, D => n2769, Z => 
                           n2767);
   U2659 : AO4 port map( A => n2549, B => n2754, C => n2635, D => n2741, Z => 
                           n2769);
   U2660 : AO4 port map( A => n2668, B => n2678, C => n2616, D => n2658, Z => 
                           n2768);
   U2661 : IV port map( A => n2602, Z => n2616);
   U2662 : AO1 port map( A => n2725, B => n2593, C => n2770, D => n2674, Z => 
                           n2766);
   U2663 : AO4 port map( A => n2771, B => n2603, C => n2645, D => n2772, Z => 
                           n2770);
   U2664 : NR2 port map( A => n2773, B => n2774, Z => n2771);
   U2665 : ND4 port map( A => n2729, B => n2775, C => n2776, D => n2777, Z => 
                           n2764);
   U2666 : ND2 port map( A => n2630, B => n2570, Z => n2777);
   U2667 : AO2 port map( A => n2778, B => n2779, C => n2725, D => n2663, Z => 
                           n2776);
   U2668 : ND2 port map( A => n2573, B => n2762, Z => n2663);
   U2669 : NR2 port map( A => n2615, B => n2644, Z => n2778);
   U2670 : ND4 port map( A => n2780, B => n2584, C => n2781, D => n2782, Z => 
                           n2775);
   U2671 : AO2 port map( A => n2688, B => n2571, C => n2612, D => n2783, Z => 
                           n2782);
   U2672 : ND3 port map( A => n2678, B => n2726, C => n2614, Z => n2781);
   U2673 : ND3 port map( A => n2661, B => n2784, C => n2594, Z => n2780);
   U2674 : AO2 port map( A => n2785, B => n2786, C => n2787, D => n2788, Z => 
                           n2763);
   U2675 : AO1 port map( A => n2561, B => n2789, C => n2790, D => n2791, Z => 
                           n2788);
   U2676 : AO6 port map( A => n2693, B => n2783, C => n2626, Z => n2791);
   U2677 : AO4 port map( A => n2558, B => n2792, C => n2607, D => n2549, Z => 
                           n2790);
   U2678 : IV port map( A => n2793, Z => n2789);
   U2679 : NR2 port map( A => n2582, B => n2636, Z => n2561);
   U2680 : AO1 port map( A => n2570, B => n2794, C => n2795, D => n2796, Z => 
                           n2787);
   U2681 : MUX21L port map( A => n2668, B => n2658, S => n2600, Z => n2795);
   U2682 : ND2 port map( A => n2797, B => n2604, Z => n2794);
   U2683 : AO1 port map( A => n2553, B => n2574, C => n2798, D => n2799, Z => 
                           n2786);
   U2684 : AO4 port map( A => n2630, B => n2603, C => n2645, D => n2800, Z => 
                           n2799);
   U2685 : AO4 port map( A => n2801, B => n2713, C => n2595, D => n2668, Z => 
                           n2798);
   U2686 : NR2 port map( A => n2698, B => n2599, Z => n2801);
   U2687 : AO1 port map( A => n2698, B => n2802, C => n2803, D => n2666, Z => 
                           n2785);
   U2688 : AO4 port map( A => n2700, B => n2626, C => n2774, D => n2558, Z => 
                           n2803);
   U2689 : IV port map( A => n2560, Z => n2700);
   U2690 : ND2 port map( A => n2669, B => n2762, Z => n2560);
   U2691 : AO3 port map( A => n2804, B => n2805, C => n2806, D => n2807, Z => 
                           n4584);
   U2692 : AO2 port map( A => n2711, B => n2808, C => n2140, D => n2107, Z => 
                           n2807);
   U2693 : AO3 port map( A => n2615, B => n2626, C => n2809, D => n2810, Z => 
                           n2808);
   U2694 : AO1 port map( A => n2811, B => n2812, C => n2813, D => n2814, Z => 
                           n2810);
   U2695 : AO6 port map( A => n2632, B => n2815, C => n2816, Z => n2814);
   U2696 : ND4 port map( A => n2625, B => n2624, C => n2817, D => n2584, Z => 
                           n2815);
   U2697 : AO4 port map( A => n2740, B => n2596, C => n2723, D => n2549, Z => 
                           n2813);
   U2698 : NR2 port map( A => n2740, B => n2774, Z => n2723);
   U2699 : OR3 port map( A => n2817, B => n2811, C => n2584, Z => n2596);
   U2700 : AO4 port map( A => n2643, B => n2668, C => n2664, D => n2603, Z => 
                           n2812);
   U2701 : EO port map( A => n2582, B => n2818, Z => n2811);
   U2702 : EO1 port map( A => n2725, B => n2635, C => n2571, D => n2645, Z => 
                           n2809);
   U2703 : ND2 port map( A => n2641, B => n2592, Z => n2571);
   U2704 : IV port map( A => n2819, Z => n2635);
   U2705 : AO2 port map( A => n2820, B => n2821, C => n2822, D => n2823, Z => 
                           n2806);
   U2706 : AO1 port map( A => n2568, B => n2574, C => n2824, D => n2825, Z => 
                           n2823);
   U2707 : IV port map( A => n2696, Z => n2825);
   U2708 : ND2 port map( A => n2750, B => n2570, Z => n2696);
   U2709 : AO1 port map( A => n2705, B => n2594, C => n2826, D => n2636, Z => 
                           n2824);
   U2710 : EON1 port map( A => n2692, B => n2592, C => n2753, D => n2688, Z => 
                           n2826);
   U2711 : ND2 port map( A => n2783, B => n2617, Z => n2574);
   U2712 : AO1 port map( A => n2599, B => n2827, C => n2674, D => n2828, Z => 
                           n2822);
   U2713 : AO6 port map( A => n2624, B => n2762, C => n2558, Z => n2828);
   U2714 : AO1 port map( A => n2829, B => n2779, C => n2830, D => n2831, Z => 
                           n2821);
   U2715 : EON1 port map( A => n2586, B => n2832, C => n2572, D => n2833, Z => 
                           n2831);
   U2716 : ND2 port map( A => n2834, B => n2584, Z => n2832);
   U2717 : EON1 port map( A => n2603, B => n2624, C => n2553, D => n2589, Z => 
                           n2830);
   U2718 : AO1 port map( A => n2568, B => n2835, C => n2836, D => n2837, Z => 
                           n2820);
   U2719 : EON1 port map( A => n2626, B => n2592, C => n2562, D => n2725, Z => 
                           n2837);
   U2720 : ND2 port map( A => n2838, B => n2546, Z => n2836);
   U2721 : IV port map( A => n2666, Z => n2546);
   U2722 : MUX21L port map( A => n2599, B => n2563, S => n2783, Z => n2838);
   U2723 : ND2 port map( A => n2644, B => n2818, Z => n2783);
   U2724 : NR4 port map( A => n2839, B => n2840, C => n2841, D => n2842, Z => 
                           n2804);
   U2725 : AO4 port map( A => n2600, B => n2668, C => n2558, D => n2640, Z => 
                           n2842);
   U2726 : EON1 port map( A => n2626, B => n2660, C => n2627, D => n2563, Z => 
                           n2841);
   U2727 : AO4 port map( A => n2819, B => n2658, C => n2549, D => n2646, Z => 
                           n2840);
   U2728 : ND2 port map( A => n2792, B => n2669, Z => n2646);
   U2729 : AO4 port map( A => n2632, B => n2800, C => n2584, D => n2843, Z => 
                           n2839);
   U2730 : ND2 port map( A => n2834, B => n2567, Z => n2843);
   U2731 : ND4 port map( A => n2844, B => n2845, C => n2846, D => n2847, Z => 
                           n4583);
   U2732 : AO1 port map( A => n2711, B => n2848, C => n2849, D => n2850, Z => 
                           n2847);
   U2733 : NR4 port map( A => n2851, B => n2852, C => n2674, D => n2675, Z => 
                           n2850);
   U2734 : AO4 port map( A => n2853, B => n2549, C => n2558, D => n2625, Z => 
                           n2675);
   U2735 : NR2 port map( A => n2774, B => n2600, Z => n2853);
   U2736 : AO4 port map( A => n2684, B => n2626, C => n2705, D => n2603, Z => 
                           n2852);
   U2737 : NR2 port map( A => n2662, B => n2589, Z => n2705);
   U2738 : AO3 port map( A => n2558, B => n2760, C => n2854, D => n2855, Z => 
                           n2851);
   U2739 : AO2 port map( A => n2615, B => n2563, C => n2553, D => n2611, Z => 
                           n2855);
   U2740 : IV port map( A => n2640, Z => n2611);
   U2741 : AO2 port map( A => n2568, B => n2856, C => n2698, D => n2772, Z => 
                           n2854);
   U2742 : ND2 port map( A => n2640, B => n2762, Z => n2772);
   U2743 : ND2 port map( A => n2835, B => n2586, Z => n2856);
   U2744 : NR2 port map( A => n4465, B => CE_I, Z => n2849);
   U2745 : ND4 port map( A => n2857, B => n2858, C => n2859, D => n2860, Z => 
                           n2848);
   U2746 : AO1 port map( A => n2736, B => n2725, C => n2861, D => n2862, Z => 
                           n2860);
   U2747 : MUX21L port map( A => n2863, B => n2864, S => n2739, Z => n2862);
   U2748 : EO port map( A => n2817, B => n2802, Z => n2739);
   U2749 : AO2 port map( A => n2568, B => n2865, C => n2599, D => n2643, Z => 
                           n2864);
   U2750 : ND2 port map( A => n2779, B => n2726, Z => n2863);
   U2751 : IV port map( A => n2605, Z => n2779);
   U2752 : AO4 port map( A => n2658, B => n2593, C => n2613, D => n2626, Z => 
                           n2861);
   U2753 : AO2 port map( A => n2653, B => n2581, C => n2563, D => n2754, Z => 
                           n2859);
   U2754 : ND2 port map( A => n2660, B => n2797, Z => n2754);
   U2755 : OR3 port map( A => n2773, B => n2829, C => n2632, Z => n2858);
   U2756 : AO7 port map( A => n2866, B => n2725, C => n2565, Z => n2857);
   U2757 : AO3 port map( A => n2867, B => n2868, C => n2619, D => n2575, Z => 
                           n2846);
   U2758 : AO4 port map( A => n2585, B => n2573, C => n2692, D => n2722, Z => 
                           n2868);
   U2759 : ND2 port map( A => n2869, B => n2745, Z => n2867);
   U2760 : ND2 port map( A => n2594, B => n2623, Z => n2745);
   U2761 : IV port map( A => n2870, Z => n2869);
   U2762 : AO6 port map( A => n2762, B => n2694, C => n2591, Z => n2870);
   U2763 : AO3 port map( A => n2793, B => n2605, C => n2871, D => n2872, Z => 
                           n2845);
   U2764 : AO6 port map( A => n2829, B => n2570, C => n2666, Z => n2872);
   U2765 : EO1 port map( A => n2873, B => n2584, C => n2694, D => n2874, Z => 
                           n2871);
   U2766 : AO6 port map( A => n2600, B => n2653, C => n2570, Z => n2874);
   U2767 : NR2 port map( A => n2584, B => n2582, Z => n2653);
   U2768 : MUX31L port map( D0 => n2875, D1 => n2819, D2 => n2724, A => n2748, 
                           B => n2876, Z => n2873);
   U2769 : NR2 port map( A => n2612, B => n2594, Z => n2876);
   U2770 : NR2 port map( A => n2589, B => n2566, Z => n2819);
   U2771 : ND2 port map( A => n2636, B => n2582, Z => n2605);
   U2772 : MUX21L port map( A => n2877, B => n2753, S => n2834, Z => n2793);
   U2773 : ND2 port map( A => n2835, B => n2617, Z => n2753);
   U2774 : ND2 port map( A => n2713, B => n2784, Z => n2877);
   U2775 : AO3 port map( A => n2878, B => n2879, C => n2636, D => n2729, Z => 
                           n2844);
   U2776 : AO4 port map( A => n2818, B => n2642, C => n2585, D => n2593, Z => 
                           n2879);
   U2777 : AO4 port map( A => n2692, B => n2722, C => n2880, D => n2591, Z => 
                           n2878);
   U2778 : AO3 port map( A => n2881, B => n2666, C => n2882, D => n2883, Z => 
                           n4582);
   U2779 : AO2 port map( A => n2629, B => n2884, C => n2140, D => n2108, Z => 
                           n2883);
   U2780 : ND4 port map( A => n2885, B => n2886, C => n2887, D => n2888, Z => 
                           n2884);
   U2781 : AO1 port map( A => n2889, B => n2599, C => n2890, D => n2891, Z => 
                           n2888);
   U2782 : NR3 port map( A => n2593, B => n2817, C => n2584, Z => n2891);
   U2783 : NR3 port map( A => n2558, B => n2590, C => n2589, Z => n2890);
   U2784 : NR2 port map( A => n2802, B => n2744, Z => n2589);
   U2785 : NR2 port map( A => n2740, B => n2736, Z => n2889);
   U2786 : IV port map( A => n2678, Z => n2736);
   U2787 : AO2 port map( A => n2630, B => n2563, C => n2662, D => n2553, Z => 
                           n2887);
   U2788 : IV port map( A => n2654, Z => n2630);
   U2789 : ND2 port map( A => n2586, B => n2694, Z => n2654);
   U2790 : AO2 port map( A => n2698, B => n2827, C => n2568, D => n2669, Z => 
                           n2886);
   U2791 : AO2 port map( A => n2721, B => n2570, C => n2716, D => n2567, Z => 
                           n2885);
   U2792 : IV port map( A => n2674, Z => n2629);
   U2793 : OR3 port map( A => n2892, B => n2680, C => n2893, Z => n2882);
   U2794 : MUX21L port map( A => n2894, B => n2895, S => n2580, Z => n2893);
   U2795 : AO3 port map( A => n2684, B => n2585, C => n2636, D => n2896, Z => 
                           n2895);
   U2796 : AO1 port map( A => n2688, B => n2717, C => n2897, D => n2898, Z => 
                           n2896);
   U2797 : AO6 port map( A => n2693, B => n2797, C => n2692, Z => n2898);
   U2798 : AN3 port map( A => n2678, B => n2624, C => n2594, Z => n2897);
   U2799 : ND2 port map( A => n2573, B => n2660, Z => n2717);
   U2800 : ND2 port map( A => n2595, B => n2802, Z => n2660);
   U2801 : NR4 port map( A => n2899, B => n2900, C => n2901, D => n2902, Z => 
                           n2894);
   U2802 : AO4 port map( A => n2744, B => n2626, C => n2623, D => n2658, Z => 
                           n2902);
   U2803 : AO6 port map( A => n2713, B => n2818, C => n2564, Z => n2623);
   U2804 : IV port map( A => n2792, Z => n2564);
   U2805 : MUX21L port map( A => n2632, B => n2645, S => n2607, Z => n2901);
   U2806 : ND2 port map( A => n2602, B => n2641, Z => n2607);
   U2807 : AO4 port map( A => n2549, B => n2573, C => n2903, D => n2603, Z => 
                           n2900);
   U2808 : AN2 port map( A => n2760, B => n2617, Z => n2903);
   U2809 : AO4 port map( A => n2558, B => n2904, C => n2668, D => n2905, Z => 
                           n2899);
   U2810 : ND2 port map( A => n2617, B => n2640, Z => n2905);
   U2811 : IV port map( A => n2662, Z => n2617);
   U2812 : NR2 port map( A => n2818, B => n2643, Z => n2662);
   U2813 : ND2 port map( A => n2678, B => n2713, Z => n2904);
   U2814 : AO1 port map( A => n2566, B => n2614, C => n2906, D => n2907, Z => 
                           n2892);
   U2815 : AO4 port map( A => n2591, B => n2800, C => n2908, D => n2692, Z => 
                           n2907);
   U2816 : NR2 port map( A => n2566, B => n2721, Z => n2908);
   U2817 : ND2 port map( A => n2722, B => n2797, Z => n2800);
   U2818 : ND2 port map( A => n2740, B => n2802, Z => n2722);
   U2819 : AO7 port map( A => n2642, B => n2726, C => n2619, Z => n2906);
   U2820 : IV port map( A => n2704, Z => n2619);
   U2821 : ND2 port map( A => n2580, B => n2584, Z => n2704);
   U2822 : NR4 port map( A => n2909, B => n2910, C => n2833, D => n2911, Z => 
                           n2881);
   U2823 : AO1 port map( A => n2626, B => n2912, C => n2740, D => n2566, Z => 
                           n2911);
   U2824 : ND2 port map( A => n2866, B => n2702, Z => n2912);
   U2825 : IV port map( A => n2797, Z => n2702);
   U2826 : ND2 port map( A => n2818, B => n2567, Z => n2797);
   U2827 : IV port map( A => n2741, Z => n2866);
   U2828 : ND2 port map( A => n2582, B => n2584, Z => n2741);
   U2829 : AO6 port map( A => n2593, B => n2760, C => n2603, Z => n2910);
   U2830 : ND2 port map( A => n2600, B => n2818, Z => n2760);
   U2831 : AO3 port map( A => n2558, B => n2573, C => n2913, D => n2914, Z => 
                           n2909);
   U2832 : MUX21L port map( A => n2563, B => n2568, S => n2915, Z => n2914);
   U2833 : AO7 port map( A => n2773, B => n2566, C => n2599, Z => n2913);
   U2834 : ND2 port map( A => n2818, B => n2865, Z => n2573);
   U2835 : AO3 port map( A => n2916, B => n2917, C => n2918, D => n2919, Z => 
                           n4581);
   U2836 : AO2 port map( A => n2711, B => n2920, C => v_SUB_WORD_0_port, D => 
                           n2140, Z => n2919);
   U2837 : ND4 port map( A => n2921, B => n2922, C => n2923, D => n2924, Z => 
                           n2920);
   U2838 : AO2 port map( A => n2925, B => n2568, C => n2915, D => n2553, Z => 
                           n2924);
   U2839 : NR2 port map( A => n2615, B => n2701, Z => n2915);
   U2840 : NR2 port map( A => n2773, B => n2829, Z => n2925);
   U2841 : IV port map( A => n2693, Z => n2829);
   U2842 : ND2 port map( A => n2643, B => n2802, Z => n2693);
   U2843 : IV port map( A => n2661, Z => n2773);
   U2844 : AO2 port map( A => n2716, B => n2926, C => n2563, D => n2669, Z => 
                           n2923);
   U2845 : ND2 port map( A => n2744, B => n2818, Z => n2669);
   U2846 : ND2 port map( A => n2792, B => n2661, Z => n2926);
   U2847 : AO2 port map( A => n2570, B => n2762, C => n2698, D => n2640, Z => 
                           n2922);
   U2848 : ND2 port map( A => n2643, B => n2818, Z => n2640);
   U2849 : ND2 port map( A => n2644, B => n2802, Z => n2762);
   U2850 : IV port map( A => n2603, Z => n2570);
   U2851 : AO2 port map( A => n2725, B => n2865, C => n2565, D => n2599, Z => 
                           n2921);
   U2852 : IV port map( A => n2549, Z => n2599);
   U2853 : IV port map( A => n2796, Z => n2711);
   U2854 : ND2 port map( A => n2575, B => n2927, Z => n2796);
   U2855 : AO2 port map( A => n2928, B => n2929, C => n2930, D => n2931, Z => 
                           n2918);
   U2856 : AO1 port map( A => n2932, B => n2678, C => n2933, D => n2833, Z => 
                           n2931);
   U2857 : NR2 port map( A => n2632, B => n2600, Z => n2833);
   U2858 : AO4 port map( A => n2549, B => n2624, C => n2591, D => n2792, Z => 
                           n2933);
   U2859 : ND2 port map( A => n2802, B => n2621, Z => n2678);
   U2860 : AO7 port map( A => n2934, B => n2692, C => n2668, Z => n2932);
   U2861 : AO1 port map( A => n2614, B => n2562, C => n2935, D => n2674, Z => 
                           n2930);
   U2862 : ND2 port map( A => n2936, B => n2580, Z => n2674);
   U2863 : AO4 port map( A => n2818, B => n2658, C => n2684, D => n2558, Z => 
                           n2935);
   U2864 : NR2 port map( A => n2565, B => n2613, Z => n2684);
   U2865 : IV port map( A => n2586, Z => n2613);
   U2866 : IV port map( A => n2624, Z => n2565);
   U2867 : ND2 port map( A => n2818, B => n2667, Z => n2624);
   U2868 : ND2 port map( A => n2694, B => n2641, Z => n2562);
   U2869 : AO1 port map( A => n2563, B => n2627, C => n2937, D => n2938, Z => 
                           n2929);
   U2870 : AO7 port map( A => n2724, B => n2668, C => n2556, Z => n2938);
   U2871 : ND2 port map( A => n2716, B => n2827, Z => n2556);
   U2872 : ND2 port map( A => n2792, B => n2694, Z => n2827);
   U2873 : ND2 port map( A => n2595, B => n2818, Z => n2694);
   U2874 : ND2 port map( A => n2664, B => n2802, Z => n2792);
   U2875 : NR2 port map( A => n2744, B => n2774, Z => n2724);
   U2876 : AO4 port map( A => n2595, B => n2658, C => n2750, D => n2549, Z => 
                           n2937);
   U2877 : NR2 port map( A => n2581, B => n2701, Z => n2750);
   U2878 : IV port map( A => n2592, Z => n2701);
   U2879 : IV port map( A => n2604, Z => n2581);
   U2880 : ND2 port map( A => n2600, B => n2802, Z => n2604);
   U2881 : IV port map( A => n2713, Z => n2600);
   U2882 : ND2 port map( A => n2625, B => n2621, Z => n2627);
   U2883 : IV port map( A => n2645, Z => n2563);
   U2884 : AO1 port map( A => n2698, B => n2875, C => n2939, D => n2666, Z => 
                           n2928);
   U2885 : ND2 port map( A => n2936, B => n2927, Z => n2666);
   U2886 : NR2 port map( A => n2940, B => n2140, Z => n2936);
   U2887 : IV port map( A => CE_I, Z => n2140);
   U2888 : AO4 port map( A => n2603, B => n2661, C => n2880, D => n2558, Z => 
                           n2939);
   U2889 : NR2 port map( A => n2567, B => n2615, Z => n2880);
   U2890 : ND2 port map( A => n2661, B => n2593, Z => n2875);
   U2891 : ND2 port map( A => n2818, B => n2726, Z => n2661);
   U2892 : AO3 port map( A => n2818, B => n2585, C => n2729, D => n2941, Z => 
                           n2917);
   U2893 : AO6 port map( A => n2816, B => n2698, C => n2942, Z => n2941);
   U2894 : AO4 port map( A => n2664, B => n2603, C => n2595, D => n2645, Z => 
                           n2942);
   U2895 : ND2 port map( A => n2614, B => n2584, Z => n2645);
   U2896 : IV port map( A => n2567, Z => n2595);
   U2897 : ND2 port map( A => n2636, B => n2614, Z => n2603);
   U2898 : IV port map( A => n2585, Z => n2614);
   U2899 : IV port map( A => n2632, Z => n2698);
   U2900 : ND2 port map( A => n2594, B => n2584, Z => n2632);
   U2901 : AO6 port map( A => n2713, B => n2818, C => n2774, Z => n2816);
   U2902 : IV port map( A => n2784, Z => n2774);
   U2903 : ND2 port map( A => n2667, B => n2802, Z => n2784);
   U2904 : IV port map( A => n2805, Z => n2729);
   U2905 : ND2 port map( A => n2575, B => n2580, Z => n2805);
   U2906 : IV port map( A => n2927, Z => n2580);
   U2907 : ND2 port map( A => n2943, B => n2944, Z => n2927);
   U2908 : AO2 port map( A => v_TEMP_VECTOR_16_port, B => n2309, C => 
                           v_TEMP_VECTOR_24_port, D => n2350, Z => n2944);
   U2909 : AO2 port map( A => v_TEMP_VECTOR_0_port, B => n2945, C => 
                           v_TEMP_VECTOR_8_port, D => n2946, Z => n2943);
   U2910 : IV port map( A => n2680, Z => n2575);
   U2911 : ND2 port map( A => CE_I, B => n2940, Z => n2680);
   U2912 : ND2 port map( A => n2947, B => n2948, Z => n2940);
   U2913 : AO2 port map( A => v_TEMP_VECTOR_22_port, B => n2309, C => 
                           v_TEMP_VECTOR_30_port, D => n2350, Z => n2948);
   U2914 : AO2 port map( A => v_TEMP_VECTOR_6_port, B => n2945, C => 
                           v_TEMP_VECTOR_14_port, D => n2946, Z => n2947);
   U2915 : ND2 port map( A => n2748, B => n2834, Z => n2585);
   U2916 : AO3 port map( A => n2549, B => n2949, C => n2950, D => n2951, Z => 
                           n2916);
   U2917 : AO2 port map( A => n2568, B => n2952, C => n2934, D => n2553, Z => 
                           n2951);
   U2918 : IV port map( A => n2658, Z => n2553);
   U2919 : ND2 port map( A => n2688, B => n2584, Z => n2658);
   U2920 : NR2 port map( A => n2590, B => n2721, Z => n2934);
   U2921 : IV port map( A => n2835, Z => n2721);
   U2922 : ND2 port map( A => n2818, B => n2664, Z => n2835);
   U2923 : IV port map( A => n2641, Z => n2590);
   U2924 : ND2 port map( A => n2744, B => n2802, Z => n2641);
   U2925 : ND2 port map( A => n2592, B => n2625, Z => n2952);
   U2926 : ND2 port map( A => n2802, B => n2567, Z => n2625);
   U2927 : ND2 port map( A => n2667, B => n2621, Z => n2567);
   U2928 : ND2 port map( A => n2818, B => n2953, Z => n2592);
   U2929 : IV port map( A => n2668, Z => n2568);
   U2930 : ND2 port map( A => n2636, B => n2612, Z => n2668);
   U2931 : AO2 port map( A => n2954, B => n2716, C => n2955, D => n2725, Z => 
                           n2950);
   U2932 : IV port map( A => n2558, Z => n2725);
   U2933 : ND2 port map( A => n2636, B => n2594, Z => n2558);
   U2934 : IV port map( A => n2642, Z => n2594);
   U2935 : ND2 port map( A => n2748, B => n2817, Z => n2642);
   U2936 : IV port map( A => n2582, Z => n2748);
   U2937 : NR2 port map( A => n2615, B => n2744, Z => n2955);
   U2938 : IV port map( A => n2621, Z => n2744);
   U2939 : ND2 port map( A => n2953, B => n2865, Z => n2621);
   U2940 : IV port map( A => n2572, Z => n2615);
   U2941 : ND2 port map( A => n2802, B => n2726, Z => n2572);
   U2942 : IV port map( A => n2626, Z => n2716);
   U2943 : ND2 port map( A => n2612, B => n2584, Z => n2626);
   U2944 : IV port map( A => n2692, Z => n2612);
   U2945 : ND2 port map( A => n2834, B => n2582, Z => n2692);
   U2946 : IV port map( A => n2817, Z => n2834);
   U2947 : NR2 port map( A => n2566, B => n2644, Z => n2954);
   U2948 : IV port map( A => n2667, Z => n2644);
   U2949 : ND2 port map( A => n2643, B => n2664, Z => n2667);
   U2950 : IV port map( A => n2593, Z => n2566);
   U2951 : ND2 port map( A => n2802, B => n2713, Z => n2593);
   U2952 : ND2 port map( A => n2664, B => n2953, Z => n2713);
   U2953 : IV port map( A => n2865, Z => n2664);
   U2954 : ND2 port map( A => n2602, B => n2586, Z => n2949);
   U2955 : ND2 port map( A => n2802, B => n2865, Z => n2586);
   U2956 : ND2 port map( A => n2740, B => n2818, Z => n2602);
   U2957 : IV port map( A => n2802, Z => n2818);
   U2958 : ND2 port map( A => n2956, B => n2957, Z => n2802);
   U2959 : AO2 port map( A => v_TEMP_VECTOR_17_port, B => n2309, C => 
                           v_TEMP_VECTOR_25_port, D => n2350, Z => n2957);
   U2960 : AO2 port map( A => v_TEMP_VECTOR_1_port, B => n2945, C => 
                           v_TEMP_VECTOR_9_port, D => n2946, Z => n2956);
   U2961 : IV port map( A => n2726, Z => n2740);
   U2962 : ND2 port map( A => n2643, B => n2865, Z => n2726);
   U2963 : ND2 port map( A => n2958, B => n2959, Z => n2865);
   U2964 : AO2 port map( A => v_TEMP_VECTOR_19_port, B => n2309, C => 
                           v_TEMP_VECTOR_27_port, D => n2350, Z => n2959);
   U2965 : AO2 port map( A => v_TEMP_VECTOR_3_port, B => n2945, C => 
                           v_TEMP_VECTOR_11_port, D => n2946, Z => n2958);
   U2966 : IV port map( A => n2953, Z => n2643);
   U2967 : ND2 port map( A => n2960, B => n2961, Z => n2953);
   U2968 : AO2 port map( A => v_TEMP_VECTOR_20_port, B => n2309, C => 
                           v_TEMP_VECTOR_28_port, D => n2350, Z => n2961);
   U2969 : AO2 port map( A => v_TEMP_VECTOR_4_port, B => n2945, C => 
                           v_TEMP_VECTOR_12_port, D => n2946, Z => n2960);
   U2970 : ND2 port map( A => n2636, B => n2688, Z => n2549);
   U2971 : IV port map( A => n2591, Z => n2688);
   U2972 : ND2 port map( A => n2582, B => n2817, Z => n2591);
   U2973 : ND2 port map( A => n2962, B => n2963, Z => n2817);
   U2974 : AO2 port map( A => v_TEMP_VECTOR_23_port, B => n2309, C => 
                           v_TEMP_VECTOR_31_port, D => n2350, Z => n2963);
   U2975 : AO2 port map( A => v_TEMP_VECTOR_7_port, B => n2945, C => 
                           v_TEMP_VECTOR_15_port, D => n2946, Z => n2962);
   U2976 : ND2 port map( A => n2964, B => n2965, Z => n2582);
   U2977 : AO2 port map( A => v_TEMP_VECTOR_18_port, B => n2309, C => 
                           v_TEMP_VECTOR_26_port, D => n2350, Z => n2965);
   U2978 : AO2 port map( A => v_TEMP_VECTOR_2_port, B => n2945, C => 
                           v_TEMP_VECTOR_10_port, D => n2946, Z => n2964);
   U2979 : IV port map( A => n2584, Z => n2636);
   U2980 : ND2 port map( A => n2966, B => n2967, Z => n2584);
   U2981 : AO2 port map( A => v_TEMP_VECTOR_21_port, B => n2309, C => 
                           v_TEMP_VECTOR_29_port, D => n2350, Z => n2967);
   U2982 : EON1 port map( A => n2137, B => n2189, C => n2537, D => n2391, Z => 
                           n2350);
   U2983 : ND2 port map( A => n2188, B => v_CALCULATION_CNTR_2_port, Z => n2137
                           );
   U2984 : IV port map( A => n2407, Z => n2188);
   U2985 : AO4 port map( A => n2397, B => n2539, C => n2398, D => n2968, Z => 
                           n2309);
   U2986 : ND2 port map( A => n2969, B => v_CALCULATION_CNTR_2_port, Z => n2968
                           );
   U2987 : AO2 port map( A => v_TEMP_VECTOR_5_port, B => n2945, C => 
                           v_TEMP_VECTOR_13_port, D => n2946, Z => n2966);
   U2988 : IV port map( A => n2261, Z => n2946);
   U2989 : AO2 port map( A => n2537, B => n2969, C => n2391, D => n2970, Z => 
                           n2261);
   U2990 : NR2 port map( A => n2407, B => v_CALCULATION_CNTR_2_port, Z => n2970
                           );
   U2991 : ND2 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n2407);
   U2992 : IV port map( A => n2189, Z => n2969);
   U2993 : AN3 port map( A => v_CALCULATION_CNTR_0_port, B => n7, C => 
                           v_CALCULATION_CNTR_2_port, Z => n2537);
   U2994 : AO4 port map( A => n2189, B => n2539, C => n2398, D => n2971, Z => 
                           n2945);
   U2995 : ND2 port map( A => n2391, B => n1036, Z => n2971);
   U2996 : IV port map( A => n2397, Z => n2391);
   U2997 : OR3 port map( A => v_CALCULATION_CNTR_4_port, B => 
                           v_CALCULATION_CNTR_3_port, C => n2540, Z => n2397);
   U2998 : ND2 port map( A => v_CALCULATION_CNTR_1_port, B => n1077, Z => n2398
                           );
   U2999 : IV port map( A => n2541, Z => n2539);
   U3000 : NR2 port map( A => n2395, B => n1036, Z => n2541);
   U3001 : ND2 port map( A => n7, B => n1077, Z => n2395);
   U3002 : OR3 port map( A => v_CALCULATION_CNTR_4_port, B => n2540, C => n1078
                           , Z => n2189);
   U3003 : OR3 port map( A => v_CALCULATION_CNTR_7_port, B => 
                           v_CALCULATION_CNTR_6_port, C => 
                           v_CALCULATION_CNTR_5_port, Z => n2540);
   U3004 : MUX21L port map( A => n4454, B => n2972, S => CE_I, Z => n4580);
   U3005 : NR2 port map( A => n2973, B => n2974, Z => n2972);
   U3006 : ND4 port map( A => n2975, B => n2976, C => n2977, D => n2978, Z => 
                           n2974);
   U3007 : NR4 port map( A => n2979, B => n2980, C => n2981, D => n2982, Z => 
                           n2978);
   U3008 : AO4 port map( A => n1080, B => n2983, C => n9, D => n2984, Z => 
                           n2982);
   U3009 : AO4 port map( A => n1081, B => n2985, C => n10, D => n2986, Z => 
                           n2981);
   U3010 : AO4 port map( A => n1082, B => n2987, C => n11, D => n2988, Z => 
                           n2980);
   U3011 : AO4 port map( A => n1083, B => n2989, C => n12, D => n2990, Z => 
                           n2979);
   U3012 : NR4 port map( A => n2991, B => n2992, C => n2993, D => n2994, Z => 
                           n2977);
   U3013 : AO4 port map( A => n1084, B => n2995, C => n13, D => n2996, Z => 
                           n2994);
   U3014 : AO4 port map( A => n1085, B => n2997, C => n14, D => n2998, Z => 
                           n2993);
   U3015 : AO4 port map( A => n1086, B => n2999, C => n15, D => n3000, Z => 
                           n2992);
   U3016 : AO4 port map( A => n1087, B => n3001, C => n16, D => n3002, Z => 
                           n2991);
   U3017 : NR4 port map( A => n3003, B => n3004, C => n3005, D => n3006, Z => 
                           n2976);
   U3018 : AO4 port map( A => n1088, B => n3007, C => n17, D => n3008, Z => 
                           n3006);
   U3019 : AO4 port map( A => n1089, B => n3009, C => n18, D => n3010, Z => 
                           n3005);
   U3020 : AO4 port map( A => n1090, B => n3011, C => n19, D => n3012, Z => 
                           n3004);
   U3021 : AO4 port map( A => n1091, B => n3013, C => n20, D => n3014, Z => 
                           n3003);
   U3022 : NR4 port map( A => n3015, B => n3016, C => n3017, D => n3018, Z => 
                           n2975);
   U3023 : AO4 port map( A => n1092, B => n3019, C => n21, D => n3020, Z => 
                           n3018);
   U3024 : AO4 port map( A => n1093, B => n3021, C => n22, D => n3022, Z => 
                           n3017);
   U3025 : AO4 port map( A => n1094, B => n3023, C => n23, D => n3024, Z => 
                           n3016);
   U3026 : AO4 port map( A => n1095, B => n3025, C => n24, D => n3026, Z => 
                           n3015);
   U3027 : ND4 port map( A => n3027, B => n3028, C => n3029, D => n3030, Z => 
                           n2973);
   U3028 : NR4 port map( A => n3031, B => n3032, C => n3033, D => n3034, Z => 
                           n3030);
   U3029 : AO4 port map( A => n1096, B => n3035, C => n25, D => n3036, Z => 
                           n3034);
   U3030 : AO4 port map( A => n1097, B => n3037, C => n26, D => n3038, Z => 
                           n3033);
   U3031 : AO4 port map( A => n1098, B => n3039, C => n27, D => n3040, Z => 
                           n3032);
   U3032 : AO4 port map( A => n1099, B => n3041, C => n28, D => n3042, Z => 
                           n3031);
   U3033 : NR4 port map( A => n3043, B => n3044, C => n3045, D => n3046, Z => 
                           n3029);
   U3034 : AO4 port map( A => n1100, B => n3047, C => n29, D => n3048, Z => 
                           n3046);
   U3035 : AO4 port map( A => n1101, B => n3049, C => n30, D => n3050, Z => 
                           n3045);
   U3036 : AO4 port map( A => n1102, B => n3051, C => n31, D => n3052, Z => 
                           n3044);
   U3037 : AO4 port map( A => n1103, B => n3053, C => n32, D => n3054, Z => 
                           n3043);
   U3038 : NR4 port map( A => n3055, B => n3056, C => n3057, D => n3058, Z => 
                           n3028);
   U3039 : AO4 port map( A => n1104, B => n3059, C => n33, D => n3060, Z => 
                           n3058);
   U3040 : AO4 port map( A => n1105, B => n3061, C => n34, D => n3062, Z => 
                           n3057);
   U3041 : AO4 port map( A => n1106, B => n3063, C => n35, D => n3064, Z => 
                           n3056);
   U3042 : AO4 port map( A => n1107, B => n3065, C => n36, D => n3066, Z => 
                           n3055);
   U3043 : NR4 port map( A => n3067, B => n3068, C => n3069, D => n3070, Z => 
                           n3027);
   U3044 : AO4 port map( A => n1108, B => n3071, C => n37, D => n3072, Z => 
                           n3070);
   U3045 : AO4 port map( A => n1109, B => n3073, C => n38, D => n3074, Z => 
                           n3069);
   U3046 : AO4 port map( A => n1110, B => n3075, C => n39, D => n3076, Z => 
                           n3068);
   U3047 : AO4 port map( A => n1111, B => n3077, C => n40, D => n3078, Z => 
                           n3067);
   U3048 : MUX21L port map( A => n1050, B => n3079, S => CE_I, Z => n4579);
   U3049 : NR2 port map( A => n3080, B => n3081, Z => n3079);
   U3050 : ND4 port map( A => n3082, B => n3083, C => n3084, D => n3085, Z => 
                           n3081);
   U3051 : NR4 port map( A => n3086, B => n3087, C => n3088, D => n3089, Z => 
                           n3085);
   U3052 : AO4 port map( A => n1112, B => n2983, C => n41, D => n2984, Z => 
                           n3089);
   U3053 : AO4 port map( A => n1113, B => n2985, C => n42, D => n2986, Z => 
                           n3088);
   U3054 : AO4 port map( A => n1114, B => n2987, C => n43, D => n2988, Z => 
                           n3087);
   U3055 : AO4 port map( A => n1115, B => n2989, C => n44, D => n2990, Z => 
                           n3086);
   U3056 : NR4 port map( A => n3090, B => n3091, C => n3092, D => n3093, Z => 
                           n3084);
   U3057 : AO4 port map( A => n1116, B => n2995, C => n45, D => n2996, Z => 
                           n3093);
   U3058 : AO4 port map( A => n1117, B => n2997, C => n46, D => n2998, Z => 
                           n3092);
   U3059 : AO4 port map( A => n1118, B => n2999, C => n47, D => n3000, Z => 
                           n3091);
   U3060 : AO4 port map( A => n1119, B => n3001, C => n48, D => n3002, Z => 
                           n3090);
   U3061 : NR4 port map( A => n3094, B => n3095, C => n3096, D => n3097, Z => 
                           n3083);
   U3062 : AO4 port map( A => n1120, B => n3007, C => n49, D => n3008, Z => 
                           n3097);
   U3063 : AO4 port map( A => n1121, B => n3009, C => n50, D => n3010, Z => 
                           n3096);
   U3064 : AO4 port map( A => n1122, B => n3011, C => n51, D => n3012, Z => 
                           n3095);
   U3065 : AO4 port map( A => n1123, B => n3013, C => n52, D => n3014, Z => 
                           n3094);
   U3066 : NR4 port map( A => n3098, B => n3099, C => n3100, D => n3101, Z => 
                           n3082);
   U3067 : AO4 port map( A => n1124, B => n3019, C => n53, D => n3020, Z => 
                           n3101);
   U3068 : AO4 port map( A => n1125, B => n3021, C => n54, D => n3022, Z => 
                           n3100);
   U3069 : AO4 port map( A => n1126, B => n3023, C => n55, D => n3024, Z => 
                           n3099);
   U3070 : AO4 port map( A => n1127, B => n3025, C => n56, D => n3026, Z => 
                           n3098);
   U3071 : ND4 port map( A => n3102, B => n3103, C => n3104, D => n3105, Z => 
                           n3080);
   U3072 : NR4 port map( A => n3106, B => n3107, C => n3108, D => n3109, Z => 
                           n3105);
   U3073 : AO4 port map( A => n1128, B => n3035, C => n57, D => n3036, Z => 
                           n3109);
   U3074 : AO4 port map( A => n1129, B => n3037, C => n58, D => n3038, Z => 
                           n3108);
   U3075 : AO4 port map( A => n1130, B => n3039, C => n59, D => n3040, Z => 
                           n3107);
   U3076 : AO4 port map( A => n1131, B => n3041, C => n60, D => n3042, Z => 
                           n3106);
   U3077 : AO4 port map( A => n3110, B => n3111, C => n3112, D => n3113, Z => 
                           n3104);
   U3078 : AO4 port map( A => n1132, B => n3047, C => n61, D => n3048, Z => 
                           n3113);
   U3079 : AO4 port map( A => n1133, B => n3049, C => n62, D => n3050, Z => 
                           n3112);
   U3080 : AO4 port map( A => n1134, B => n3051, C => n63, D => n3052, Z => 
                           n3111);
   U3081 : AO4 port map( A => n1135, B => n3053, C => n64, D => n3054, Z => 
                           n3110);
   U3082 : NR4 port map( A => n3114, B => n3115, C => n3116, D => n3117, Z => 
                           n3103);
   U3083 : AO4 port map( A => n1136, B => n3059, C => n65, D => n3060, Z => 
                           n3117);
   U3084 : AO4 port map( A => n1137, B => n3061, C => n66, D => n3062, Z => 
                           n3116);
   U3085 : AO4 port map( A => n1138, B => n3063, C => n67, D => n3064, Z => 
                           n3115);
   U3086 : AO4 port map( A => n1139, B => n3065, C => n68, D => n3066, Z => 
                           n3114);
   U3087 : NR4 port map( A => n3118, B => n3119, C => n3120, D => n3121, Z => 
                           n3102);
   U3088 : AO4 port map( A => n1140, B => n3071, C => n69, D => n3072, Z => 
                           n3121);
   U3089 : AO4 port map( A => n1141, B => n3073, C => n70, D => n3074, Z => 
                           n3120);
   U3090 : AO4 port map( A => n1142, B => n3075, C => n71, D => n3076, Z => 
                           n3119);
   U3091 : AO4 port map( A => n1143, B => n3077, C => n72, D => n3078, Z => 
                           n3118);
   U3092 : MUX21L port map( A => n1059, B => n3122, S => CE_I, Z => n4578);
   U3093 : NR2 port map( A => n3123, B => n3124, Z => n3122);
   U3094 : ND4 port map( A => n3125, B => n3126, C => n3127, D => n3128, Z => 
                           n3124);
   U3095 : NR4 port map( A => n3129, B => n3130, C => n3131, D => n3132, Z => 
                           n3128);
   U3096 : AO4 port map( A => n1144, B => n2983, C => n73, D => n2984, Z => 
                           n3132);
   U3097 : AO4 port map( A => n1145, B => n2985, C => n74, D => n2986, Z => 
                           n3131);
   U3098 : AO4 port map( A => n1146, B => n2987, C => n75, D => n2988, Z => 
                           n3130);
   U3099 : AO4 port map( A => n1147, B => n2989, C => n76, D => n2990, Z => 
                           n3129);
   U3100 : NR4 port map( A => n3133, B => n3134, C => n3135, D => n3136, Z => 
                           n3127);
   U3101 : AO4 port map( A => n1148, B => n2995, C => n77, D => n2996, Z => 
                           n3136);
   U3102 : AO4 port map( A => n1149, B => n2997, C => n78, D => n2998, Z => 
                           n3135);
   U3103 : AO4 port map( A => n1150, B => n2999, C => n79, D => n3000, Z => 
                           n3134);
   U3104 : AO4 port map( A => n1151, B => n3001, C => n80, D => n3002, Z => 
                           n3133);
   U3105 : NR4 port map( A => n3137, B => n3138, C => n3139, D => n3140, Z => 
                           n3126);
   U3106 : AO4 port map( A => n1152, B => n3007, C => n81, D => n3008, Z => 
                           n3140);
   U3107 : AO4 port map( A => n1153, B => n3009, C => n82, D => n3010, Z => 
                           n3139);
   U3108 : AO4 port map( A => n1154, B => n3011, C => n83, D => n3012, Z => 
                           n3138);
   U3109 : AO4 port map( A => n1155, B => n3013, C => n84, D => n3014, Z => 
                           n3137);
   U3110 : NR4 port map( A => n3141, B => n3142, C => n3143, D => n3144, Z => 
                           n3125);
   U3111 : AO4 port map( A => n1156, B => n3019, C => n85, D => n3020, Z => 
                           n3144);
   U3112 : AO4 port map( A => n1157, B => n3021, C => n86, D => n3022, Z => 
                           n3143);
   U3113 : AO4 port map( A => n1158, B => n3023, C => n87, D => n3024, Z => 
                           n3142);
   U3114 : AO4 port map( A => n1159, B => n3025, C => n88, D => n3026, Z => 
                           n3141);
   U3115 : ND4 port map( A => n3145, B => n3146, C => n3147, D => n3148, Z => 
                           n3123);
   U3116 : NR4 port map( A => n3149, B => n3150, C => n3151, D => n3152, Z => 
                           n3148);
   U3117 : AO4 port map( A => n1160, B => n3035, C => n89, D => n3036, Z => 
                           n3152);
   U3118 : AO4 port map( A => n1161, B => n3037, C => n90, D => n3038, Z => 
                           n3151);
   U3119 : AO4 port map( A => n1162, B => n3039, C => n91, D => n3040, Z => 
                           n3150);
   U3120 : AO4 port map( A => n1163, B => n3041, C => n92, D => n3042, Z => 
                           n3149);
   U3121 : NR4 port map( A => n3153, B => n3154, C => n3155, D => n3156, Z => 
                           n3147);
   U3122 : AO4 port map( A => n1164, B => n3047, C => n93, D => n3048, Z => 
                           n3156);
   U3123 : AO4 port map( A => n1165, B => n3049, C => n94, D => n3050, Z => 
                           n3155);
   U3124 : AO4 port map( A => n1166, B => n3051, C => n95, D => n3052, Z => 
                           n3154);
   U3125 : AO4 port map( A => n1167, B => n3053, C => n96, D => n3054, Z => 
                           n3153);
   U3126 : NR4 port map( A => n3157, B => n3158, C => n3159, D => n3160, Z => 
                           n3146);
   U3127 : AO4 port map( A => n1168, B => n3059, C => n97, D => n3060, Z => 
                           n3160);
   U3128 : AO4 port map( A => n1169, B => n3061, C => n98, D => n3062, Z => 
                           n3159);
   U3129 : AO4 port map( A => n1170, B => n3063, C => n99, D => n3064, Z => 
                           n3158);
   U3130 : AO4 port map( A => n1171, B => n3065, C => n100, D => n3066, Z => 
                           n3157);
   U3131 : NR4 port map( A => n3161, B => n3162, C => n3163, D => n3164, Z => 
                           n3145);
   U3132 : AO4 port map( A => n1172, B => n3071, C => n101, D => n3072, Z => 
                           n3164);
   U3133 : AO4 port map( A => n1173, B => n3073, C => n102, D => n3074, Z => 
                           n3163);
   U3134 : AO4 port map( A => n1174, B => n3075, C => n103, D => n3076, Z => 
                           n3162);
   U3135 : AO4 port map( A => n1175, B => n3077, C => n104, D => n3078, Z => 
                           n3161);
   U3136 : MUX21L port map( A => n1068, B => n3165, S => CE_I, Z => n4577);
   U3137 : NR2 port map( A => n3166, B => n3167, Z => n3165);
   U3138 : ND4 port map( A => n3168, B => n3169, C => n3170, D => n3171, Z => 
                           n3167);
   U3139 : NR4 port map( A => n3172, B => n3173, C => n3174, D => n3175, Z => 
                           n3171);
   U3140 : AO4 port map( A => n1176, B => n2983, C => n105, D => n2984, Z => 
                           n3175);
   U3141 : AO4 port map( A => n1177, B => n2985, C => n106, D => n2986, Z => 
                           n3174);
   U3142 : AO4 port map( A => n1178, B => n2987, C => n107, D => n2988, Z => 
                           n3173);
   U3143 : AO4 port map( A => n1179, B => n2989, C => n108, D => n2990, Z => 
                           n3172);
   U3144 : NR4 port map( A => n3176, B => n3177, C => n3178, D => n3179, Z => 
                           n3170);
   U3145 : AO4 port map( A => n1180, B => n2995, C => n109, D => n2996, Z => 
                           n3179);
   U3146 : AO4 port map( A => n1181, B => n2997, C => n110, D => n2998, Z => 
                           n3178);
   U3147 : AO4 port map( A => n1182, B => n2999, C => n111, D => n3000, Z => 
                           n3177);
   U3148 : AO4 port map( A => n1183, B => n3001, C => n112, D => n3002, Z => 
                           n3176);
   U3149 : NR4 port map( A => n3180, B => n3181, C => n3182, D => n3183, Z => 
                           n3169);
   U3150 : AO4 port map( A => n1184, B => n3007, C => n113, D => n3008, Z => 
                           n3183);
   U3151 : AO4 port map( A => n1185, B => n3009, C => n114, D => n3010, Z => 
                           n3182);
   U3152 : AO4 port map( A => n1186, B => n3011, C => n115, D => n3012, Z => 
                           n3181);
   U3153 : AO4 port map( A => n1187, B => n3013, C => n116, D => n3014, Z => 
                           n3180);
   U3154 : NR4 port map( A => n3184, B => n3185, C => n3186, D => n3187, Z => 
                           n3168);
   U3155 : AO4 port map( A => n1188, B => n3019, C => n117, D => n3020, Z => 
                           n3187);
   U3156 : AO4 port map( A => n1189, B => n3021, C => n118, D => n3022, Z => 
                           n3186);
   U3157 : AO4 port map( A => n1190, B => n3023, C => n119, D => n3024, Z => 
                           n3185);
   U3158 : AO4 port map( A => n1191, B => n3025, C => n120, D => n3026, Z => 
                           n3184);
   U3159 : ND4 port map( A => n3188, B => n3189, C => n3190, D => n3191, Z => 
                           n3166);
   U3160 : NR4 port map( A => n3192, B => n3193, C => n3194, D => n3195, Z => 
                           n3191);
   U3161 : AO4 port map( A => n1192, B => n3035, C => n121, D => n3036, Z => 
                           n3195);
   U3162 : AO4 port map( A => n1193, B => n3037, C => n122, D => n3038, Z => 
                           n3194);
   U3163 : AO4 port map( A => n1194, B => n3039, C => n123, D => n3040, Z => 
                           n3193);
   U3164 : AO4 port map( A => n1195, B => n3041, C => n124, D => n3042, Z => 
                           n3192);
   U3165 : NR4 port map( A => n3196, B => n3197, C => n3198, D => n3199, Z => 
                           n3190);
   U3166 : AO4 port map( A => n1196, B => n3047, C => n125, D => n3048, Z => 
                           n3199);
   U3167 : AO4 port map( A => n1197, B => n3049, C => n126, D => n3050, Z => 
                           n3198);
   U3168 : AO4 port map( A => n1198, B => n3051, C => n127, D => n3052, Z => 
                           n3197);
   U3169 : AO4 port map( A => n1199, B => n3053, C => n128, D => n3054, Z => 
                           n3196);
   U3170 : NR4 port map( A => n3200, B => n3201, C => n3202, D => n3203, Z => 
                           n3189);
   U3171 : AO4 port map( A => n1200, B => n3059, C => n129, D => n3060, Z => 
                           n3203);
   U3172 : AO4 port map( A => n1201, B => n3061, C => n130, D => n3062, Z => 
                           n3202);
   U3173 : AO4 port map( A => n1202, B => n3063, C => n131, D => n3064, Z => 
                           n3201);
   U3174 : AO4 port map( A => n1203, B => n3065, C => n132, D => n3066, Z => 
                           n3200);
   U3175 : NR4 port map( A => n3204, B => n3205, C => n3206, D => n3207, Z => 
                           n3188);
   U3176 : AO4 port map( A => n1204, B => n3071, C => n133, D => n3072, Z => 
                           n3207);
   U3177 : AO4 port map( A => n1205, B => n3073, C => n134, D => n3074, Z => 
                           n3206);
   U3178 : AO4 port map( A => n1206, B => n3075, C => n135, D => n3076, Z => 
                           n3205);
   U3179 : AO4 port map( A => n1207, B => n3077, C => n136, D => n3078, Z => 
                           n3204);
   U3180 : MUX21L port map( A => n4457, B => n3208, S => CE_I, Z => n4576);
   U3181 : NR2 port map( A => n3209, B => n3210, Z => n3208);
   U3182 : ND4 port map( A => n3211, B => n3212, C => n3213, D => n3214, Z => 
                           n3210);
   U3183 : NR4 port map( A => n3215, B => n3216, C => n3217, D => n3218, Z => 
                           n3214);
   U3184 : AO4 port map( A => n1208, B => n2983, C => n137, D => n2984, Z => 
                           n3218);
   U3185 : AO4 port map( A => n1209, B => n2985, C => n138, D => n2986, Z => 
                           n3217);
   U3186 : AO4 port map( A => n1210, B => n2987, C => n139, D => n2988, Z => 
                           n3216);
   U3187 : AO4 port map( A => n1211, B => n2989, C => n140, D => n2990, Z => 
                           n3215);
   U3188 : NR4 port map( A => n3219, B => n3220, C => n3221, D => n3222, Z => 
                           n3213);
   U3189 : AO4 port map( A => n1212, B => n2995, C => n141, D => n2996, Z => 
                           n3222);
   U3190 : AO4 port map( A => n1213, B => n2997, C => n142, D => n2998, Z => 
                           n3221);
   U3191 : AO4 port map( A => n1214, B => n2999, C => n143, D => n3000, Z => 
                           n3220);
   U3192 : AO4 port map( A => n1215, B => n3001, C => n144, D => n3002, Z => 
                           n3219);
   U3193 : NR4 port map( A => n3223, B => n3224, C => n3225, D => n3226, Z => 
                           n3212);
   U3194 : AO4 port map( A => n1216, B => n3007, C => n145, D => n3008, Z => 
                           n3226);
   U3195 : AO4 port map( A => n1217, B => n3009, C => n146, D => n3010, Z => 
                           n3225);
   U3196 : AO4 port map( A => n1218, B => n3011, C => n147, D => n3012, Z => 
                           n3224);
   U3197 : AO4 port map( A => n1219, B => n3013, C => n148, D => n3014, Z => 
                           n3223);
   U3198 : NR4 port map( A => n3227, B => n3228, C => n3229, D => n3230, Z => 
                           n3211);
   U3199 : AO4 port map( A => n1220, B => n3019, C => n149, D => n3020, Z => 
                           n3230);
   U3200 : AO4 port map( A => n1221, B => n3021, C => n150, D => n3022, Z => 
                           n3229);
   U3201 : AO4 port map( A => n1222, B => n3023, C => n151, D => n3024, Z => 
                           n3228);
   U3202 : AO4 port map( A => n1223, B => n3025, C => n152, D => n3026, Z => 
                           n3227);
   U3203 : ND4 port map( A => n3231, B => n3232, C => n3233, D => n3234, Z => 
                           n3209);
   U3204 : NR4 port map( A => n3235, B => n3236, C => n3237, D => n3238, Z => 
                           n3234);
   U3205 : AO4 port map( A => n1224, B => n3035, C => n153, D => n3036, Z => 
                           n3238);
   U3206 : AO4 port map( A => n1225, B => n3037, C => n154, D => n3038, Z => 
                           n3237);
   U3207 : AO4 port map( A => n1226, B => n3039, C => n155, D => n3040, Z => 
                           n3236);
   U3208 : AO4 port map( A => n1227, B => n3041, C => n156, D => n3042, Z => 
                           n3235);
   U3209 : NR4 port map( A => n3239, B => n3240, C => n3241, D => n3242, Z => 
                           n3233);
   U3210 : AO4 port map( A => n1228, B => n3047, C => n157, D => n3048, Z => 
                           n3242);
   U3211 : AO4 port map( A => n1229, B => n3049, C => n158, D => n3050, Z => 
                           n3241);
   U3212 : AO4 port map( A => n1230, B => n3051, C => n159, D => n3052, Z => 
                           n3240);
   U3213 : AO4 port map( A => n1231, B => n3053, C => n160, D => n3054, Z => 
                           n3239);
   U3214 : NR4 port map( A => n3243, B => n3244, C => n3245, D => n3246, Z => 
                           n3232);
   U3215 : AO4 port map( A => n1232, B => n3059, C => n161, D => n3060, Z => 
                           n3246);
   U3216 : AO4 port map( A => n1233, B => n3061, C => n162, D => n3062, Z => 
                           n3245);
   U3217 : AO4 port map( A => n1234, B => n3063, C => n163, D => n3064, Z => 
                           n3244);
   U3218 : AO4 port map( A => n1235, B => n3065, C => n164, D => n3066, Z => 
                           n3243);
   U3219 : NR4 port map( A => n3247, B => n3248, C => n3249, D => n3250, Z => 
                           n3231);
   U3220 : AO4 port map( A => n1236, B => n3071, C => n165, D => n3072, Z => 
                           n3250);
   U3221 : AO4 port map( A => n1237, B => n3073, C => n166, D => n3074, Z => 
                           n3249);
   U3222 : AO4 port map( A => n1238, B => n3075, C => n167, D => n3076, Z => 
                           n3248);
   U3223 : AO4 port map( A => n1239, B => n3077, C => n168, D => n3078, Z => 
                           n3247);
   U3224 : MUX21L port map( A => n1051, B => n3251, S => CE_I, Z => n4575);
   U3225 : NR2 port map( A => n3252, B => n3253, Z => n3251);
   U3226 : ND4 port map( A => n3254, B => n3255, C => n3256, D => n3257, Z => 
                           n3253);
   U3227 : NR4 port map( A => n3258, B => n3259, C => n3260, D => n3261, Z => 
                           n3257);
   U3228 : AO4 port map( A => n1240, B => n2983, C => n169, D => n2984, Z => 
                           n3261);
   U3229 : AO4 port map( A => n1241, B => n2985, C => n170, D => n2986, Z => 
                           n3260);
   U3230 : AO4 port map( A => n1242, B => n2987, C => n171, D => n2988, Z => 
                           n3259);
   U3231 : AO4 port map( A => n1243, B => n2989, C => n172, D => n2990, Z => 
                           n3258);
   U3232 : NR4 port map( A => n3262, B => n3263, C => n3264, D => n3265, Z => 
                           n3256);
   U3233 : AO4 port map( A => n1244, B => n2995, C => n173, D => n2996, Z => 
                           n3265);
   U3234 : AO4 port map( A => n1245, B => n2997, C => n174, D => n2998, Z => 
                           n3264);
   U3235 : AO4 port map( A => n1246, B => n2999, C => n175, D => n3000, Z => 
                           n3263);
   U3236 : AO4 port map( A => n1247, B => n3001, C => n176, D => n3002, Z => 
                           n3262);
   U3237 : NR4 port map( A => n3266, B => n3267, C => n3268, D => n3269, Z => 
                           n3255);
   U3238 : AO4 port map( A => n1248, B => n3007, C => n177, D => n3008, Z => 
                           n3269);
   U3239 : AO4 port map( A => n1249, B => n3009, C => n178, D => n3010, Z => 
                           n3268);
   U3240 : AO4 port map( A => n1250, B => n3011, C => n179, D => n3012, Z => 
                           n3267);
   U3241 : AO4 port map( A => n1251, B => n3013, C => n180, D => n3014, Z => 
                           n3266);
   U3242 : NR4 port map( A => n3270, B => n3271, C => n3272, D => n3273, Z => 
                           n3254);
   U3243 : AO4 port map( A => n1252, B => n3019, C => n181, D => n3020, Z => 
                           n3273);
   U3244 : AO4 port map( A => n1253, B => n3021, C => n182, D => n3022, Z => 
                           n3272);
   U3245 : AO4 port map( A => n1254, B => n3023, C => n183, D => n3024, Z => 
                           n3271);
   U3246 : AO4 port map( A => n1255, B => n3025, C => n184, D => n3026, Z => 
                           n3270);
   U3247 : ND4 port map( A => n3274, B => n3275, C => n3276, D => n3277, Z => 
                           n3252);
   U3248 : NR4 port map( A => n3278, B => n3279, C => n3280, D => n3281, Z => 
                           n3277);
   U3249 : AO4 port map( A => n1256, B => n3035, C => n185, D => n3036, Z => 
                           n3281);
   U3250 : AO4 port map( A => n1257, B => n3037, C => n186, D => n3038, Z => 
                           n3280);
   U3251 : AO4 port map( A => n1258, B => n3039, C => n187, D => n3040, Z => 
                           n3279);
   U3252 : AO4 port map( A => n1259, B => n3041, C => n188, D => n3042, Z => 
                           n3278);
   U3253 : NR4 port map( A => n3282, B => n3283, C => n3284, D => n3285, Z => 
                           n3276);
   U3254 : AO4 port map( A => n1260, B => n3047, C => n189, D => n3048, Z => 
                           n3285);
   U3255 : AO4 port map( A => n1261, B => n3049, C => n190, D => n3050, Z => 
                           n3284);
   U3256 : AO4 port map( A => n1262, B => n3051, C => n191, D => n3052, Z => 
                           n3283);
   U3257 : AO4 port map( A => n1263, B => n3053, C => n192, D => n3054, Z => 
                           n3282);
   U3258 : NR4 port map( A => n3286, B => n3287, C => n3288, D => n3289, Z => 
                           n3275);
   U3259 : AO4 port map( A => n1264, B => n3059, C => n193, D => n3060, Z => 
                           n3289);
   U3260 : AO4 port map( A => n1265, B => n3061, C => n194, D => n3062, Z => 
                           n3288);
   U3261 : AO4 port map( A => n1266, B => n3063, C => n195, D => n3064, Z => 
                           n3287);
   U3262 : AO4 port map( A => n1267, B => n3065, C => n196, D => n3066, Z => 
                           n3286);
   U3263 : NR4 port map( A => n3290, B => n3291, C => n3292, D => n3293, Z => 
                           n3274);
   U3264 : AO4 port map( A => n1268, B => n3071, C => n197, D => n3072, Z => 
                           n3293);
   U3265 : AO4 port map( A => n1269, B => n3073, C => n198, D => n3074, Z => 
                           n3292);
   U3266 : AO4 port map( A => n1270, B => n3075, C => n199, D => n3076, Z => 
                           n3291);
   U3267 : AO4 port map( A => n1271, B => n3077, C => n200, D => n3078, Z => 
                           n3290);
   U3268 : MUX21L port map( A => n1060, B => n3294, S => CE_I, Z => n4574);
   U3269 : NR2 port map( A => n3295, B => n3296, Z => n3294);
   U3270 : ND4 port map( A => n3297, B => n3298, C => n3299, D => n3300, Z => 
                           n3296);
   U3271 : NR4 port map( A => n3301, B => n3302, C => n3303, D => n3304, Z => 
                           n3300);
   U3272 : AO4 port map( A => n1272, B => n2983, C => n201, D => n2984, Z => 
                           n3304);
   U3273 : AO4 port map( A => n1273, B => n2985, C => n202, D => n2986, Z => 
                           n3303);
   U3274 : AO4 port map( A => n1274, B => n2987, C => n203, D => n2988, Z => 
                           n3302);
   U3275 : AO4 port map( A => n1275, B => n2989, C => n204, D => n2990, Z => 
                           n3301);
   U3276 : NR4 port map( A => n3305, B => n3306, C => n3307, D => n3308, Z => 
                           n3299);
   U3277 : AO4 port map( A => n1276, B => n2995, C => n205, D => n2996, Z => 
                           n3308);
   U3278 : AO4 port map( A => n1277, B => n2997, C => n206, D => n2998, Z => 
                           n3307);
   U3279 : AO4 port map( A => n1278, B => n2999, C => n207, D => n3000, Z => 
                           n3306);
   U3280 : AO4 port map( A => n1279, B => n3001, C => n208, D => n3002, Z => 
                           n3305);
   U3281 : NR4 port map( A => n3309, B => n3310, C => n3311, D => n3312, Z => 
                           n3298);
   U3282 : AO4 port map( A => n1280, B => n3007, C => n209, D => n3008, Z => 
                           n3312);
   U3283 : AO4 port map( A => n1281, B => n3009, C => n210, D => n3010, Z => 
                           n3311);
   U3284 : AO4 port map( A => n1282, B => n3011, C => n211, D => n3012, Z => 
                           n3310);
   U3285 : AO4 port map( A => n1283, B => n3013, C => n212, D => n3014, Z => 
                           n3309);
   U3286 : NR4 port map( A => n3313, B => n3314, C => n3315, D => n3316, Z => 
                           n3297);
   U3287 : AO4 port map( A => n1284, B => n3019, C => n213, D => n3020, Z => 
                           n3316);
   U3288 : AO4 port map( A => n1285, B => n3021, C => n214, D => n3022, Z => 
                           n3315);
   U3289 : AO4 port map( A => n1286, B => n3023, C => n215, D => n3024, Z => 
                           n3314);
   U3290 : AO4 port map( A => n1287, B => n3025, C => n216, D => n3026, Z => 
                           n3313);
   U3291 : ND4 port map( A => n3317, B => n3318, C => n3319, D => n3320, Z => 
                           n3295);
   U3292 : NR4 port map( A => n3321, B => n3322, C => n3323, D => n3324, Z => 
                           n3320);
   U3293 : AO4 port map( A => n1288, B => n3035, C => n217, D => n3036, Z => 
                           n3324);
   U3294 : AO4 port map( A => n1289, B => n3037, C => n218, D => n3038, Z => 
                           n3323);
   U3295 : AO4 port map( A => n1290, B => n3039, C => n219, D => n3040, Z => 
                           n3322);
   U3296 : AO4 port map( A => n1291, B => n3041, C => n220, D => n3042, Z => 
                           n3321);
   U3297 : NR4 port map( A => n3325, B => n3326, C => n3327, D => n3328, Z => 
                           n3319);
   U3298 : AO4 port map( A => n1292, B => n3047, C => n221, D => n3048, Z => 
                           n3328);
   U3299 : AO4 port map( A => n1293, B => n3049, C => n222, D => n3050, Z => 
                           n3327);
   U3300 : AO4 port map( A => n1294, B => n3051, C => n223, D => n3052, Z => 
                           n3326);
   U3301 : AO4 port map( A => n1295, B => n3053, C => n224, D => n3054, Z => 
                           n3325);
   U3302 : NR4 port map( A => n3329, B => n3330, C => n3331, D => n3332, Z => 
                           n3318);
   U3303 : AO4 port map( A => n1296, B => n3059, C => n225, D => n3060, Z => 
                           n3332);
   U3304 : AO4 port map( A => n1297, B => n3061, C => n226, D => n3062, Z => 
                           n3331);
   U3305 : AO4 port map( A => n1298, B => n3063, C => n227, D => n3064, Z => 
                           n3330);
   U3306 : AO4 port map( A => n1299, B => n3065, C => n228, D => n3066, Z => 
                           n3329);
   U3307 : NR4 port map( A => n3333, B => n3334, C => n3335, D => n3336, Z => 
                           n3317);
   U3308 : AO4 port map( A => n1300, B => n3071, C => n229, D => n3072, Z => 
                           n3336);
   U3309 : AO4 port map( A => n1301, B => n3073, C => n230, D => n3074, Z => 
                           n3335);
   U3310 : AO4 port map( A => n1302, B => n3075, C => n231, D => n3076, Z => 
                           n3334);
   U3311 : AO4 port map( A => n1303, B => n3077, C => n232, D => n3078, Z => 
                           n3333);
   U3312 : MUX21L port map( A => n1069, B => n3337, S => CE_I, Z => n4573);
   U3313 : NR2 port map( A => n3338, B => n3339, Z => n3337);
   U3314 : ND4 port map( A => n3340, B => n3341, C => n3342, D => n3343, Z => 
                           n3339);
   U3315 : NR4 port map( A => n3344, B => n3345, C => n3346, D => n3347, Z => 
                           n3343);
   U3316 : AO4 port map( A => n1304, B => n2983, C => n233, D => n2984, Z => 
                           n3347);
   U3317 : AO4 port map( A => n1305, B => n2985, C => n234, D => n2986, Z => 
                           n3346);
   U3318 : AO4 port map( A => n1306, B => n2987, C => n235, D => n2988, Z => 
                           n3345);
   U3319 : AO4 port map( A => n1307, B => n2989, C => n236, D => n2990, Z => 
                           n3344);
   U3320 : NR4 port map( A => n3348, B => n3349, C => n3350, D => n3351, Z => 
                           n3342);
   U3321 : AO4 port map( A => n1308, B => n2995, C => n237, D => n2996, Z => 
                           n3351);
   U3322 : AO4 port map( A => n1309, B => n2997, C => n238, D => n2998, Z => 
                           n3350);
   U3323 : AO4 port map( A => n1310, B => n2999, C => n239, D => n3000, Z => 
                           n3349);
   U3324 : AO4 port map( A => n1311, B => n3001, C => n240, D => n3002, Z => 
                           n3348);
   U3325 : NR4 port map( A => n3352, B => n3353, C => n3354, D => n3355, Z => 
                           n3341);
   U3326 : AO4 port map( A => n1312, B => n3007, C => n241, D => n3008, Z => 
                           n3355);
   U3327 : AO4 port map( A => n1313, B => n3009, C => n242, D => n3010, Z => 
                           n3354);
   U3328 : AO4 port map( A => n1314, B => n3011, C => n243, D => n3012, Z => 
                           n3353);
   U3329 : AO4 port map( A => n1315, B => n3013, C => n244, D => n3014, Z => 
                           n3352);
   U3330 : NR4 port map( A => n3356, B => n3357, C => n3358, D => n3359, Z => 
                           n3340);
   U3331 : AO4 port map( A => n1316, B => n3019, C => n245, D => n3020, Z => 
                           n3359);
   U3332 : AO4 port map( A => n1317, B => n3021, C => n246, D => n3022, Z => 
                           n3358);
   U3333 : AO4 port map( A => n1318, B => n3023, C => n247, D => n3024, Z => 
                           n3357);
   U3334 : AO4 port map( A => n1319, B => n3025, C => n248, D => n3026, Z => 
                           n3356);
   U3335 : ND4 port map( A => n3360, B => n3361, C => n3362, D => n3363, Z => 
                           n3338);
   U3336 : NR4 port map( A => n3364, B => n3365, C => n3366, D => n3367, Z => 
                           n3363);
   U3337 : AO4 port map( A => n1320, B => n3035, C => n249, D => n3036, Z => 
                           n3367);
   U3338 : AO4 port map( A => n1321, B => n3037, C => n250, D => n3038, Z => 
                           n3366);
   U3339 : AO4 port map( A => n1322, B => n3039, C => n251, D => n3040, Z => 
                           n3365);
   U3340 : AO4 port map( A => n1323, B => n3041, C => n252, D => n3042, Z => 
                           n3364);
   U3341 : NR4 port map( A => n3368, B => n3369, C => n3370, D => n3371, Z => 
                           n3362);
   U3342 : AO4 port map( A => n1324, B => n3047, C => n253, D => n3048, Z => 
                           n3371);
   U3343 : AO4 port map( A => n1325, B => n3049, C => n254, D => n3050, Z => 
                           n3370);
   U3344 : AO4 port map( A => n1326, B => n3051, C => n255, D => n3052, Z => 
                           n3369);
   U3345 : AO4 port map( A => n1327, B => n3053, C => n256, D => n3054, Z => 
                           n3368);
   U3346 : NR4 port map( A => n3372, B => n3373, C => n3374, D => n3375, Z => 
                           n3361);
   U3347 : AO4 port map( A => n1328, B => n3059, C => n257, D => n3060, Z => 
                           n3375);
   U3348 : AO4 port map( A => n1329, B => n3061, C => n258, D => n3062, Z => 
                           n3374);
   U3349 : AO4 port map( A => n1330, B => n3063, C => n259, D => n3064, Z => 
                           n3373);
   U3350 : AO4 port map( A => n1331, B => n3065, C => n260, D => n3066, Z => 
                           n3372);
   U3351 : NR4 port map( A => n3376, B => n3377, C => n3378, D => n3379, Z => 
                           n3360);
   U3352 : AO4 port map( A => n1332, B => n3071, C => n261, D => n3072, Z => 
                           n3379);
   U3353 : AO4 port map( A => n1333, B => n3073, C => n262, D => n3074, Z => 
                           n3378);
   U3354 : AO4 port map( A => n1334, B => n3075, C => n263, D => n3076, Z => 
                           n3377);
   U3355 : AO4 port map( A => n1335, B => n3077, C => n264, D => n3078, Z => 
                           n3376);
   U3356 : MUX21L port map( A => n1047, B => n3380, S => CE_I, Z => n4572);
   U3357 : NR2 port map( A => n3381, B => n3382, Z => n3380);
   U3358 : ND4 port map( A => n3383, B => n3384, C => n3385, D => n3386, Z => 
                           n3382);
   U3359 : NR4 port map( A => n3387, B => n3388, C => n3389, D => n3390, Z => 
                           n3386);
   U3360 : AO4 port map( A => n1336, B => n2983, C => n265, D => n2984, Z => 
                           n3390);
   U3361 : AO4 port map( A => n1337, B => n2985, C => n266, D => n2986, Z => 
                           n3389);
   U3362 : AO4 port map( A => n1338, B => n2987, C => n267, D => n2988, Z => 
                           n3388);
   U3363 : AO4 port map( A => n1339, B => n2989, C => n268, D => n2990, Z => 
                           n3387);
   U3364 : NR4 port map( A => n3391, B => n3392, C => n3393, D => n3394, Z => 
                           n3385);
   U3365 : AO4 port map( A => n1340, B => n2995, C => n269, D => n2996, Z => 
                           n3394);
   U3366 : AO4 port map( A => n1341, B => n2997, C => n270, D => n2998, Z => 
                           n3393);
   U3367 : AO4 port map( A => n1342, B => n2999, C => n271, D => n3000, Z => 
                           n3392);
   U3368 : AO4 port map( A => n1343, B => n3001, C => n272, D => n3002, Z => 
                           n3391);
   U3369 : NR4 port map( A => n3395, B => n3396, C => n3397, D => n3398, Z => 
                           n3384);
   U3370 : AO4 port map( A => n1344, B => n3007, C => n273, D => n3008, Z => 
                           n3398);
   U3371 : AO4 port map( A => n1345, B => n3009, C => n274, D => n3010, Z => 
                           n3397);
   U3372 : AO4 port map( A => n1346, B => n3011, C => n275, D => n3012, Z => 
                           n3396);
   U3373 : AO4 port map( A => n1347, B => n3013, C => n276, D => n3014, Z => 
                           n3395);
   U3374 : NR4 port map( A => n3399, B => n3400, C => n3401, D => n3402, Z => 
                           n3383);
   U3375 : AO4 port map( A => n1348, B => n3019, C => n277, D => n3020, Z => 
                           n3402);
   U3376 : AO4 port map( A => n1349, B => n3021, C => n278, D => n3022, Z => 
                           n3401);
   U3377 : AO4 port map( A => n1350, B => n3023, C => n279, D => n3024, Z => 
                           n3400);
   U3378 : AO4 port map( A => n1351, B => n3025, C => n280, D => n3026, Z => 
                           n3399);
   U3379 : ND4 port map( A => n3403, B => n3404, C => n3405, D => n3406, Z => 
                           n3381);
   U3380 : NR4 port map( A => n3407, B => n3408, C => n3409, D => n3410, Z => 
                           n3406);
   U3381 : AO4 port map( A => n1352, B => n3035, C => n281, D => n3036, Z => 
                           n3410);
   U3382 : AO4 port map( A => n1353, B => n3037, C => n282, D => n3038, Z => 
                           n3409);
   U3383 : AO4 port map( A => n1354, B => n3039, C => n283, D => n3040, Z => 
                           n3408);
   U3384 : AO4 port map( A => n1355, B => n3041, C => n284, D => n3042, Z => 
                           n3407);
   U3385 : NR4 port map( A => n3411, B => n3412, C => n3413, D => n3414, Z => 
                           n3405);
   U3386 : AO4 port map( A => n1356, B => n3047, C => n285, D => n3048, Z => 
                           n3414);
   U3387 : AO4 port map( A => n1357, B => n3049, C => n286, D => n3050, Z => 
                           n3413);
   U3388 : AO4 port map( A => n1358, B => n3051, C => n287, D => n3052, Z => 
                           n3412);
   U3389 : AO4 port map( A => n1359, B => n3053, C => n288, D => n3054, Z => 
                           n3411);
   U3390 : NR4 port map( A => n3415, B => n3416, C => n3417, D => n3418, Z => 
                           n3404);
   U3391 : AO4 port map( A => n1360, B => n3059, C => n289, D => n3060, Z => 
                           n3418);
   U3392 : AO4 port map( A => n1361, B => n3061, C => n290, D => n3062, Z => 
                           n3417);
   U3393 : AO4 port map( A => n1362, B => n3063, C => n291, D => n3064, Z => 
                           n3416);
   U3394 : AO4 port map( A => n1363, B => n3065, C => n292, D => n3066, Z => 
                           n3415);
   U3395 : NR4 port map( A => n3419, B => n3420, C => n3421, D => n3422, Z => 
                           n3403);
   U3396 : AO4 port map( A => n1364, B => n3071, C => n293, D => n3072, Z => 
                           n3422);
   U3397 : AO4 port map( A => n1365, B => n3073, C => n294, D => n3074, Z => 
                           n3421);
   U3398 : AO4 port map( A => n1366, B => n3075, C => n295, D => n3076, Z => 
                           n3420);
   U3399 : AO4 port map( A => n1367, B => n3077, C => n296, D => n3078, Z => 
                           n3419);
   U3400 : MUX21L port map( A => n1053, B => n3423, S => CE_I, Z => n4571);
   U3401 : NR2 port map( A => n3424, B => n3425, Z => n3423);
   U3402 : ND4 port map( A => n3426, B => n3427, C => n3428, D => n3429, Z => 
                           n3425);
   U3403 : NR4 port map( A => n3430, B => n3431, C => n3432, D => n3433, Z => 
                           n3429);
   U3404 : AO4 port map( A => n1368, B => n2983, C => n297, D => n2984, Z => 
                           n3433);
   U3405 : AO4 port map( A => n1369, B => n2985, C => n298, D => n2986, Z => 
                           n3432);
   U3406 : AO4 port map( A => n1370, B => n2987, C => n299, D => n2988, Z => 
                           n3431);
   U3407 : AO4 port map( A => n1371, B => n2989, C => n300, D => n2990, Z => 
                           n3430);
   U3408 : NR4 port map( A => n3434, B => n3435, C => n3436, D => n3437, Z => 
                           n3428);
   U3409 : AO4 port map( A => n1372, B => n2995, C => n301, D => n2996, Z => 
                           n3437);
   U3410 : AO4 port map( A => n1373, B => n2997, C => n302, D => n2998, Z => 
                           n3436);
   U3411 : AO4 port map( A => n1374, B => n2999, C => n303, D => n3000, Z => 
                           n3435);
   U3412 : AO4 port map( A => n1375, B => n3001, C => n304, D => n3002, Z => 
                           n3434);
   U3413 : NR4 port map( A => n3438, B => n3439, C => n3440, D => n3441, Z => 
                           n3427);
   U3414 : AO4 port map( A => n1376, B => n3007, C => n305, D => n3008, Z => 
                           n3441);
   U3415 : AO4 port map( A => n1377, B => n3009, C => n306, D => n3010, Z => 
                           n3440);
   U3416 : AO4 port map( A => n1378, B => n3011, C => n307, D => n3012, Z => 
                           n3439);
   U3417 : AO4 port map( A => n1379, B => n3013, C => n308, D => n3014, Z => 
                           n3438);
   U3418 : NR4 port map( A => n3442, B => n3443, C => n3444, D => n3445, Z => 
                           n3426);
   U3419 : AO4 port map( A => n1380, B => n3019, C => n309, D => n3020, Z => 
                           n3445);
   U3420 : AO4 port map( A => n1381, B => n3021, C => n310, D => n3022, Z => 
                           n3444);
   U3421 : AO4 port map( A => n1382, B => n3023, C => n311, D => n3024, Z => 
                           n3443);
   U3422 : AO4 port map( A => n1383, B => n3025, C => n312, D => n3026, Z => 
                           n3442);
   U3423 : ND4 port map( A => n3446, B => n3447, C => n3448, D => n3449, Z => 
                           n3424);
   U3424 : NR4 port map( A => n3450, B => n3451, C => n3452, D => n3453, Z => 
                           n3449);
   U3425 : AO4 port map( A => n1384, B => n3035, C => n313, D => n3036, Z => 
                           n3453);
   U3426 : AO4 port map( A => n1385, B => n3037, C => n314, D => n3038, Z => 
                           n3452);
   U3427 : AO4 port map( A => n1386, B => n3039, C => n315, D => n3040, Z => 
                           n3451);
   U3428 : AO4 port map( A => n1387, B => n3041, C => n316, D => n3042, Z => 
                           n3450);
   U3429 : NR4 port map( A => n3454, B => n3455, C => n3456, D => n3457, Z => 
                           n3448);
   U3430 : AO4 port map( A => n1388, B => n3047, C => n317, D => n3048, Z => 
                           n3457);
   U3431 : AO4 port map( A => n1389, B => n3049, C => n318, D => n3050, Z => 
                           n3456);
   U3432 : AO4 port map( A => n1390, B => n3051, C => n319, D => n3052, Z => 
                           n3455);
   U3433 : AO4 port map( A => n1391, B => n3053, C => n320, D => n3054, Z => 
                           n3454);
   U3434 : NR4 port map( A => n3458, B => n3459, C => n3460, D => n3461, Z => 
                           n3447);
   U3435 : AO4 port map( A => n1392, B => n3059, C => n321, D => n3060, Z => 
                           n3461);
   U3436 : AO4 port map( A => n1393, B => n3061, C => n322, D => n3062, Z => 
                           n3460);
   U3437 : AO4 port map( A => n1394, B => n3063, C => n323, D => n3064, Z => 
                           n3459);
   U3438 : AO4 port map( A => n1395, B => n3065, C => n324, D => n3066, Z => 
                           n3458);
   U3439 : NR4 port map( A => n3462, B => n3463, C => n3464, D => n3465, Z => 
                           n3446);
   U3440 : AO4 port map( A => n1396, B => n3071, C => n325, D => n3072, Z => 
                           n3465);
   U3441 : AO4 port map( A => n1397, B => n3073, C => n326, D => n3074, Z => 
                           n3464);
   U3442 : AO4 port map( A => n1398, B => n3075, C => n327, D => n3076, Z => 
                           n3463);
   U3443 : AO4 port map( A => n1399, B => n3077, C => n328, D => n3078, Z => 
                           n3462);
   U3444 : MUX21L port map( A => n1061, B => n3466, S => CE_I, Z => n4570);
   U3445 : NR2 port map( A => n3467, B => n3468, Z => n3466);
   U3446 : ND4 port map( A => n3469, B => n3470, C => n3471, D => n3472, Z => 
                           n3468);
   U3447 : NR4 port map( A => n3473, B => n3474, C => n3475, D => n3476, Z => 
                           n3472);
   U3448 : AO4 port map( A => n1400, B => n2983, C => n329, D => n2984, Z => 
                           n3476);
   U3449 : AO4 port map( A => n1401, B => n2985, C => n330, D => n2986, Z => 
                           n3475);
   U3450 : AO4 port map( A => n1402, B => n2987, C => n331, D => n2988, Z => 
                           n3474);
   U3451 : AO4 port map( A => n1403, B => n2989, C => n332, D => n2990, Z => 
                           n3473);
   U3452 : NR4 port map( A => n3477, B => n3478, C => n3479, D => n3480, Z => 
                           n3471);
   U3453 : AO4 port map( A => n1404, B => n2995, C => n333, D => n2996, Z => 
                           n3480);
   U3454 : AO4 port map( A => n1405, B => n2997, C => n334, D => n2998, Z => 
                           n3479);
   U3455 : AO4 port map( A => n1406, B => n2999, C => n335, D => n3000, Z => 
                           n3478);
   U3456 : AO4 port map( A => n1407, B => n3001, C => n336, D => n3002, Z => 
                           n3477);
   U3457 : NR4 port map( A => n3481, B => n3482, C => n3483, D => n3484, Z => 
                           n3470);
   U3458 : AO4 port map( A => n1408, B => n3007, C => n337, D => n3008, Z => 
                           n3484);
   U3459 : AO4 port map( A => n1409, B => n3009, C => n338, D => n3010, Z => 
                           n3483);
   U3460 : AO4 port map( A => n1410, B => n3011, C => n339, D => n3012, Z => 
                           n3482);
   U3461 : AO4 port map( A => n1411, B => n3013, C => n340, D => n3014, Z => 
                           n3481);
   U3462 : NR4 port map( A => n3485, B => n3486, C => n3487, D => n3488, Z => 
                           n3469);
   U3463 : AO4 port map( A => n1412, B => n3019, C => n341, D => n3020, Z => 
                           n3488);
   U3464 : AO4 port map( A => n1413, B => n3021, C => n342, D => n3022, Z => 
                           n3487);
   U3465 : AO4 port map( A => n1414, B => n3023, C => n343, D => n3024, Z => 
                           n3486);
   U3466 : AO4 port map( A => n1415, B => n3025, C => n344, D => n3026, Z => 
                           n3485);
   U3467 : ND4 port map( A => n3489, B => n3490, C => n3491, D => n3492, Z => 
                           n3467);
   U3468 : NR4 port map( A => n3493, B => n3494, C => n3495, D => n3496, Z => 
                           n3492);
   U3469 : AO4 port map( A => n1416, B => n3035, C => n345, D => n3036, Z => 
                           n3496);
   U3470 : AO4 port map( A => n1417, B => n3037, C => n346, D => n3038, Z => 
                           n3495);
   U3471 : AO4 port map( A => n1418, B => n3039, C => n347, D => n3040, Z => 
                           n3494);
   U3472 : AO4 port map( A => n1419, B => n3041, C => n348, D => n3042, Z => 
                           n3493);
   U3473 : NR4 port map( A => n3497, B => n3498, C => n3499, D => n3500, Z => 
                           n3491);
   U3474 : AO4 port map( A => n1420, B => n3047, C => n349, D => n3048, Z => 
                           n3500);
   U3475 : AO4 port map( A => n1421, B => n3049, C => n350, D => n3050, Z => 
                           n3499);
   U3476 : AO4 port map( A => n1422, B => n3051, C => n351, D => n3052, Z => 
                           n3498);
   U3477 : AO4 port map( A => n1423, B => n3053, C => n352, D => n3054, Z => 
                           n3497);
   U3478 : NR4 port map( A => n3501, B => n3502, C => n3503, D => n3504, Z => 
                           n3490);
   U3479 : AO4 port map( A => n1424, B => n3059, C => n353, D => n3060, Z => 
                           n3504);
   U3480 : AO4 port map( A => n1425, B => n3061, C => n354, D => n3062, Z => 
                           n3503);
   U3481 : AO4 port map( A => n1426, B => n3063, C => n355, D => n3064, Z => 
                           n3502);
   U3482 : AO4 port map( A => n1427, B => n3065, C => n356, D => n3066, Z => 
                           n3501);
   U3483 : NR4 port map( A => n3505, B => n3506, C => n3507, D => n3508, Z => 
                           n3489);
   U3484 : AO4 port map( A => n1428, B => n3071, C => n357, D => n3072, Z => 
                           n3508);
   U3485 : AO4 port map( A => n1429, B => n3073, C => n358, D => n3074, Z => 
                           n3507);
   U3486 : AO4 port map( A => n1430, B => n3075, C => n359, D => n3076, Z => 
                           n3506);
   U3487 : AO4 port map( A => n1431, B => n3077, C => n360, D => n3078, Z => 
                           n3505);
   U3488 : MUX21L port map( A => n1070, B => n3509, S => CE_I, Z => n4569);
   U3489 : NR2 port map( A => n3510, B => n3511, Z => n3509);
   U3490 : ND4 port map( A => n3512, B => n3513, C => n3514, D => n3515, Z => 
                           n3511);
   U3491 : NR4 port map( A => n3516, B => n3517, C => n3518, D => n3519, Z => 
                           n3515);
   U3492 : AO4 port map( A => n1432, B => n2983, C => n361, D => n2984, Z => 
                           n3519);
   U3493 : AO4 port map( A => n1433, B => n2985, C => n362, D => n2986, Z => 
                           n3518);
   U3494 : AO4 port map( A => n1434, B => n2987, C => n363, D => n2988, Z => 
                           n3517);
   U3495 : AO4 port map( A => n1435, B => n2989, C => n364, D => n2990, Z => 
                           n3516);
   U3496 : NR4 port map( A => n3520, B => n3521, C => n3522, D => n3523, Z => 
                           n3514);
   U3497 : AO4 port map( A => n1436, B => n2995, C => n365, D => n2996, Z => 
                           n3523);
   U3498 : AO4 port map( A => n1437, B => n2997, C => n366, D => n2998, Z => 
                           n3522);
   U3499 : AO4 port map( A => n1438, B => n2999, C => n367, D => n3000, Z => 
                           n3521);
   U3500 : AO4 port map( A => n1439, B => n3001, C => n368, D => n3002, Z => 
                           n3520);
   U3501 : NR4 port map( A => n3524, B => n3525, C => n3526, D => n3527, Z => 
                           n3513);
   U3502 : AO4 port map( A => n1440, B => n3007, C => n369, D => n3008, Z => 
                           n3527);
   U3503 : AO4 port map( A => n1441, B => n3009, C => n370, D => n3010, Z => 
                           n3526);
   U3504 : AO4 port map( A => n1442, B => n3011, C => n371, D => n3012, Z => 
                           n3525);
   U3505 : AO4 port map( A => n1443, B => n3013, C => n372, D => n3014, Z => 
                           n3524);
   U3506 : NR4 port map( A => n3528, B => n3529, C => n3530, D => n3531, Z => 
                           n3512);
   U3507 : AO4 port map( A => n1444, B => n3019, C => n373, D => n3020, Z => 
                           n3531);
   U3508 : AO4 port map( A => n1445, B => n3021, C => n374, D => n3022, Z => 
                           n3530);
   U3509 : AO4 port map( A => n1446, B => n3023, C => n375, D => n3024, Z => 
                           n3529);
   U3510 : AO4 port map( A => n1447, B => n3025, C => n376, D => n3026, Z => 
                           n3528);
   U3511 : ND4 port map( A => n3532, B => n3533, C => n3534, D => n3535, Z => 
                           n3510);
   U3512 : NR4 port map( A => n3536, B => n3537, C => n3538, D => n3539, Z => 
                           n3535);
   U3513 : AO4 port map( A => n1448, B => n3035, C => n377, D => n3036, Z => 
                           n3539);
   U3514 : AO4 port map( A => n1449, B => n3037, C => n378, D => n3038, Z => 
                           n3538);
   U3515 : AO4 port map( A => n1450, B => n3039, C => n379, D => n3040, Z => 
                           n3537);
   U3516 : AO4 port map( A => n1451, B => n3041, C => n380, D => n3042, Z => 
                           n3536);
   U3517 : NR4 port map( A => n3540, B => n3541, C => n3542, D => n3543, Z => 
                           n3534);
   U3518 : AO4 port map( A => n1452, B => n3047, C => n381, D => n3048, Z => 
                           n3543);
   U3519 : AO4 port map( A => n1453, B => n3049, C => n382, D => n3050, Z => 
                           n3542);
   U3520 : AO4 port map( A => n1454, B => n3051, C => n383, D => n3052, Z => 
                           n3541);
   U3521 : AO4 port map( A => n1455, B => n3053, C => n384, D => n3054, Z => 
                           n3540);
   U3522 : NR4 port map( A => n3544, B => n3545, C => n3546, D => n3547, Z => 
                           n3533);
   U3523 : AO4 port map( A => n1456, B => n3059, C => n385, D => n3060, Z => 
                           n3547);
   U3524 : AO4 port map( A => n1457, B => n3061, C => n386, D => n3062, Z => 
                           n3546);
   U3525 : AO4 port map( A => n1458, B => n3063, C => n387, D => n3064, Z => 
                           n3545);
   U3526 : AO4 port map( A => n1459, B => n3065, C => n388, D => n3066, Z => 
                           n3544);
   U3527 : NR4 port map( A => n3548, B => n3549, C => n3550, D => n3551, Z => 
                           n3532);
   U3528 : AO4 port map( A => n1460, B => n3071, C => n389, D => n3072, Z => 
                           n3551);
   U3529 : AO4 port map( A => n1461, B => n3073, C => n390, D => n3074, Z => 
                           n3550);
   U3530 : AO4 port map( A => n1462, B => n3075, C => n391, D => n3076, Z => 
                           n3549);
   U3531 : AO4 port map( A => n1463, B => n3077, C => n392, D => n3078, Z => 
                           n3548);
   U3532 : MUX21L port map( A => n1048, B => n3552, S => CE_I, Z => n4568);
   U3533 : NR2 port map( A => n3553, B => n3554, Z => n3552);
   U3534 : ND4 port map( A => n3555, B => n3556, C => n3557, D => n3558, Z => 
                           n3554);
   U3535 : NR4 port map( A => n3559, B => n3560, C => n3561, D => n3562, Z => 
                           n3558);
   U3536 : AO4 port map( A => n1464, B => n2983, C => n393, D => n2984, Z => 
                           n3562);
   U3537 : AO4 port map( A => n1465, B => n2985, C => n394, D => n2986, Z => 
                           n3561);
   U3538 : AO4 port map( A => n1466, B => n2987, C => n395, D => n2988, Z => 
                           n3560);
   U3539 : AO4 port map( A => n1467, B => n2989, C => n396, D => n2990, Z => 
                           n3559);
   U3540 : NR4 port map( A => n3563, B => n3564, C => n3565, D => n3566, Z => 
                           n3557);
   U3541 : AO4 port map( A => n1468, B => n2995, C => n397, D => n2996, Z => 
                           n3566);
   U3542 : AO4 port map( A => n1469, B => n2997, C => n398, D => n2998, Z => 
                           n3565);
   U3543 : AO4 port map( A => n1470, B => n2999, C => n399, D => n3000, Z => 
                           n3564);
   U3544 : AO4 port map( A => n1471, B => n3001, C => n400, D => n3002, Z => 
                           n3563);
   U3545 : NR4 port map( A => n3567, B => n3568, C => n3569, D => n3570, Z => 
                           n3556);
   U3546 : AO4 port map( A => n1472, B => n3007, C => n401, D => n3008, Z => 
                           n3570);
   U3547 : AO4 port map( A => n1473, B => n3009, C => n402, D => n3010, Z => 
                           n3569);
   U3548 : AO4 port map( A => n1474, B => n3011, C => n403, D => n3012, Z => 
                           n3568);
   U3549 : AO4 port map( A => n1475, B => n3013, C => n404, D => n3014, Z => 
                           n3567);
   U3550 : NR4 port map( A => n3571, B => n3572, C => n3573, D => n3574, Z => 
                           n3555);
   U3551 : AO4 port map( A => n1476, B => n3019, C => n405, D => n3020, Z => 
                           n3574);
   U3552 : AO4 port map( A => n1477, B => n3021, C => n406, D => n3022, Z => 
                           n3573);
   U3553 : AO4 port map( A => n1478, B => n3023, C => n407, D => n3024, Z => 
                           n3572);
   U3554 : AO4 port map( A => n1479, B => n3025, C => n408, D => n3026, Z => 
                           n3571);
   U3555 : ND4 port map( A => n3575, B => n3576, C => n3577, D => n3578, Z => 
                           n3553);
   U3556 : NR4 port map( A => n3579, B => n3580, C => n3581, D => n3582, Z => 
                           n3578);
   U3557 : AO4 port map( A => n1480, B => n3035, C => n409, D => n3036, Z => 
                           n3582);
   U3558 : AO4 port map( A => n1481, B => n3037, C => n410, D => n3038, Z => 
                           n3581);
   U3559 : AO4 port map( A => n1482, B => n3039, C => n411, D => n3040, Z => 
                           n3580);
   U3560 : AO4 port map( A => n1483, B => n3041, C => n412, D => n3042, Z => 
                           n3579);
   U3561 : NR4 port map( A => n3583, B => n3584, C => n3585, D => n3586, Z => 
                           n3577);
   U3562 : AO4 port map( A => n1484, B => n3047, C => n413, D => n3048, Z => 
                           n3586);
   U3563 : AO4 port map( A => n1485, B => n3049, C => n414, D => n3050, Z => 
                           n3585);
   U3564 : AO4 port map( A => n1486, B => n3051, C => n415, D => n3052, Z => 
                           n3584);
   U3565 : AO4 port map( A => n1487, B => n3053, C => n416, D => n3054, Z => 
                           n3583);
   U3566 : NR4 port map( A => n3587, B => n3588, C => n3589, D => n3590, Z => 
                           n3576);
   U3567 : AO4 port map( A => n1488, B => n3059, C => n417, D => n3060, Z => 
                           n3590);
   U3568 : AO4 port map( A => n1489, B => n3061, C => n418, D => n3062, Z => 
                           n3589);
   U3569 : AO4 port map( A => n1490, B => n3063, C => n419, D => n3064, Z => 
                           n3588);
   U3570 : AO4 port map( A => n1491, B => n3065, C => n420, D => n3066, Z => 
                           n3587);
   U3571 : NR4 port map( A => n3591, B => n3592, C => n3593, D => n3594, Z => 
                           n3575);
   U3572 : AO4 port map( A => n1492, B => n3071, C => n421, D => n3072, Z => 
                           n3594);
   U3573 : AO4 port map( A => n1493, B => n3073, C => n422, D => n3074, Z => 
                           n3593);
   U3574 : AO4 port map( A => n1494, B => n3075, C => n423, D => n3076, Z => 
                           n3592);
   U3575 : AO4 port map( A => n1495, B => n3077, C => n424, D => n3078, Z => 
                           n3591);
   U3576 : MUX21L port map( A => n1054, B => n3595, S => CE_I, Z => n4567);
   U3577 : NR2 port map( A => n3596, B => n3597, Z => n3595);
   U3578 : ND4 port map( A => n3598, B => n3599, C => n3600, D => n3601, Z => 
                           n3597);
   U3579 : NR4 port map( A => n3602, B => n3603, C => n3604, D => n3605, Z => 
                           n3601);
   U3580 : AO4 port map( A => n1496, B => n2983, C => n425, D => n2984, Z => 
                           n3605);
   U3581 : AO4 port map( A => n1497, B => n2985, C => n426, D => n2986, Z => 
                           n3604);
   U3582 : AO4 port map( A => n1498, B => n2987, C => n427, D => n2988, Z => 
                           n3603);
   U3583 : AO4 port map( A => n1499, B => n2989, C => n428, D => n2990, Z => 
                           n3602);
   U3584 : NR4 port map( A => n3606, B => n3607, C => n3608, D => n3609, Z => 
                           n3600);
   U3585 : AO4 port map( A => n1500, B => n2995, C => n429, D => n2996, Z => 
                           n3609);
   U3586 : AO4 port map( A => n1501, B => n2997, C => n430, D => n2998, Z => 
                           n3608);
   U3587 : AO4 port map( A => n1502, B => n2999, C => n431, D => n3000, Z => 
                           n3607);
   U3588 : AO4 port map( A => n1503, B => n3001, C => n432, D => n3002, Z => 
                           n3606);
   U3589 : NR4 port map( A => n3610, B => n3611, C => n3612, D => n3613, Z => 
                           n3599);
   U3590 : AO4 port map( A => n1504, B => n3007, C => n433, D => n3008, Z => 
                           n3613);
   U3591 : AO4 port map( A => n1505, B => n3009, C => n434, D => n3010, Z => 
                           n3612);
   U3592 : AO4 port map( A => n1506, B => n3011, C => n435, D => n3012, Z => 
                           n3611);
   U3593 : AO4 port map( A => n1507, B => n3013, C => n436, D => n3014, Z => 
                           n3610);
   U3594 : NR4 port map( A => n3614, B => n3615, C => n3616, D => n3617, Z => 
                           n3598);
   U3595 : AO4 port map( A => n1508, B => n3019, C => n437, D => n3020, Z => 
                           n3617);
   U3596 : AO4 port map( A => n1509, B => n3021, C => n438, D => n3022, Z => 
                           n3616);
   U3597 : AO4 port map( A => n1510, B => n3023, C => n439, D => n3024, Z => 
                           n3615);
   U3598 : AO4 port map( A => n1511, B => n3025, C => n440, D => n3026, Z => 
                           n3614);
   U3599 : ND4 port map( A => n3618, B => n3619, C => n3620, D => n3621, Z => 
                           n3596);
   U3600 : NR4 port map( A => n3622, B => n3623, C => n3624, D => n3625, Z => 
                           n3621);
   U3601 : AO4 port map( A => n1512, B => n3035, C => n441, D => n3036, Z => 
                           n3625);
   U3602 : AO4 port map( A => n1513, B => n3037, C => n442, D => n3038, Z => 
                           n3624);
   U3603 : AO4 port map( A => n1514, B => n3039, C => n443, D => n3040, Z => 
                           n3623);
   U3604 : AO4 port map( A => n1515, B => n3041, C => n444, D => n3042, Z => 
                           n3622);
   U3605 : NR4 port map( A => n3626, B => n3627, C => n3628, D => n3629, Z => 
                           n3620);
   U3606 : AO4 port map( A => n1516, B => n3047, C => n445, D => n3048, Z => 
                           n3629);
   U3607 : AO4 port map( A => n1517, B => n3049, C => n446, D => n3050, Z => 
                           n3628);
   U3608 : AO4 port map( A => n1518, B => n3051, C => n447, D => n3052, Z => 
                           n3627);
   U3609 : AO4 port map( A => n1519, B => n3053, C => n448, D => n3054, Z => 
                           n3626);
   U3610 : NR4 port map( A => n3630, B => n3631, C => n3632, D => n3633, Z => 
                           n3619);
   U3611 : AO4 port map( A => n1520, B => n3059, C => n449, D => n3060, Z => 
                           n3633);
   U3612 : AO4 port map( A => n1521, B => n3061, C => n450, D => n3062, Z => 
                           n3632);
   U3613 : AO4 port map( A => n1522, B => n3063, C => n451, D => n3064, Z => 
                           n3631);
   U3614 : AO4 port map( A => n1523, B => n3065, C => n452, D => n3066, Z => 
                           n3630);
   U3615 : NR4 port map( A => n3634, B => n3635, C => n3636, D => n3637, Z => 
                           n3618);
   U3616 : AO4 port map( A => n1524, B => n3071, C => n453, D => n3072, Z => 
                           n3637);
   U3617 : AO4 port map( A => n1525, B => n3073, C => n454, D => n3074, Z => 
                           n3636);
   U3618 : AO4 port map( A => n1526, B => n3075, C => n455, D => n3076, Z => 
                           n3635);
   U3619 : AO4 port map( A => n1527, B => n3077, C => n456, D => n3078, Z => 
                           n3634);
   U3620 : MUX21L port map( A => n1062, B => n3638, S => CE_I, Z => n4566);
   U3621 : NR2 port map( A => n3639, B => n3640, Z => n3638);
   U3622 : ND4 port map( A => n3641, B => n3642, C => n3643, D => n3644, Z => 
                           n3640);
   U3623 : NR4 port map( A => n3645, B => n3646, C => n3647, D => n3648, Z => 
                           n3644);
   U3624 : AO4 port map( A => n1528, B => n2983, C => n457, D => n2984, Z => 
                           n3648);
   U3625 : AO4 port map( A => n1529, B => n2985, C => n458, D => n2986, Z => 
                           n3647);
   U3626 : AO4 port map( A => n1530, B => n2987, C => n459, D => n2988, Z => 
                           n3646);
   U3627 : AO4 port map( A => n1531, B => n2989, C => n460, D => n2990, Z => 
                           n3645);
   U3628 : NR4 port map( A => n3649, B => n3650, C => n3651, D => n3652, Z => 
                           n3643);
   U3629 : AO4 port map( A => n1532, B => n2995, C => n461, D => n2996, Z => 
                           n3652);
   U3630 : AO4 port map( A => n1533, B => n2997, C => n462, D => n2998, Z => 
                           n3651);
   U3631 : AO4 port map( A => n1534, B => n2999, C => n463, D => n3000, Z => 
                           n3650);
   U3632 : AO4 port map( A => n1535, B => n3001, C => n464, D => n3002, Z => 
                           n3649);
   U3633 : NR4 port map( A => n3653, B => n3654, C => n3655, D => n3656, Z => 
                           n3642);
   U3634 : AO4 port map( A => n1536, B => n3007, C => n465, D => n3008, Z => 
                           n3656);
   U3635 : AO4 port map( A => n1537, B => n3009, C => n466, D => n3010, Z => 
                           n3655);
   U3636 : AO4 port map( A => n1538, B => n3011, C => n467, D => n3012, Z => 
                           n3654);
   U3637 : AO4 port map( A => n1539, B => n3013, C => n468, D => n3014, Z => 
                           n3653);
   U3638 : NR4 port map( A => n3657, B => n3658, C => n3659, D => n3660, Z => 
                           n3641);
   U3639 : AO4 port map( A => n1540, B => n3019, C => n469, D => n3020, Z => 
                           n3660);
   U3640 : AO4 port map( A => n1541, B => n3021, C => n470, D => n3022, Z => 
                           n3659);
   U3641 : AO4 port map( A => n1542, B => n3023, C => n471, D => n3024, Z => 
                           n3658);
   U3642 : AO4 port map( A => n1543, B => n3025, C => n472, D => n3026, Z => 
                           n3657);
   U3643 : ND4 port map( A => n3661, B => n3662, C => n3663, D => n3664, Z => 
                           n3639);
   U3644 : NR4 port map( A => n3665, B => n3666, C => n3667, D => n3668, Z => 
                           n3664);
   U3645 : AO4 port map( A => n1544, B => n3035, C => n473, D => n3036, Z => 
                           n3668);
   U3646 : AO4 port map( A => n1545, B => n3037, C => n474, D => n3038, Z => 
                           n3667);
   U3647 : AO4 port map( A => n1546, B => n3039, C => n475, D => n3040, Z => 
                           n3666);
   U3648 : AO4 port map( A => n1547, B => n3041, C => n476, D => n3042, Z => 
                           n3665);
   U3649 : NR4 port map( A => n3669, B => n3670, C => n3671, D => n3672, Z => 
                           n3663);
   U3650 : AO4 port map( A => n1548, B => n3047, C => n477, D => n3048, Z => 
                           n3672);
   U3651 : AO4 port map( A => n1549, B => n3049, C => n478, D => n3050, Z => 
                           n3671);
   U3652 : AO4 port map( A => n1550, B => n3051, C => n479, D => n3052, Z => 
                           n3670);
   U3653 : AO4 port map( A => n1551, B => n3053, C => n480, D => n3054, Z => 
                           n3669);
   U3654 : NR4 port map( A => n3673, B => n3674, C => n3675, D => n3676, Z => 
                           n3662);
   U3655 : AO4 port map( A => n1552, B => n3059, C => n481, D => n3060, Z => 
                           n3676);
   U3656 : AO4 port map( A => n1553, B => n3061, C => n482, D => n3062, Z => 
                           n3675);
   U3657 : AO4 port map( A => n1554, B => n3063, C => n483, D => n3064, Z => 
                           n3674);
   U3658 : AO4 port map( A => n1555, B => n3065, C => n484, D => n3066, Z => 
                           n3673);
   U3659 : NR4 port map( A => n3677, B => n3678, C => n3679, D => n3680, Z => 
                           n3661);
   U3660 : AO4 port map( A => n1556, B => n3071, C => n485, D => n3072, Z => 
                           n3680);
   U3661 : AO4 port map( A => n1557, B => n3073, C => n486, D => n3074, Z => 
                           n3679);
   U3662 : AO4 port map( A => n1558, B => n3075, C => n487, D => n3076, Z => 
                           n3678);
   U3663 : AO4 port map( A => n1559, B => n3077, C => n488, D => n3078, Z => 
                           n3677);
   U3664 : MUX21L port map( A => n1071, B => n3681, S => CE_I, Z => n4565);
   U3665 : NR2 port map( A => n3682, B => n3683, Z => n3681);
   U3666 : ND4 port map( A => n3684, B => n3685, C => n3686, D => n3687, Z => 
                           n3683);
   U3667 : NR4 port map( A => n3688, B => n3689, C => n3690, D => n3691, Z => 
                           n3687);
   U3668 : AO4 port map( A => n1560, B => n2983, C => n489, D => n2984, Z => 
                           n3691);
   U3669 : AO4 port map( A => n1561, B => n2985, C => n490, D => n2986, Z => 
                           n3690);
   U3670 : AO4 port map( A => n1562, B => n2987, C => n491, D => n2988, Z => 
                           n3689);
   U3671 : AO4 port map( A => n1563, B => n2989, C => n492, D => n2990, Z => 
                           n3688);
   U3672 : NR4 port map( A => n3692, B => n3693, C => n3694, D => n3695, Z => 
                           n3686);
   U3673 : AO4 port map( A => n1564, B => n2995, C => n493, D => n2996, Z => 
                           n3695);
   U3674 : AO4 port map( A => n1565, B => n2997, C => n494, D => n2998, Z => 
                           n3694);
   U3675 : AO4 port map( A => n1566, B => n2999, C => n495, D => n3000, Z => 
                           n3693);
   U3676 : AO4 port map( A => n1567, B => n3001, C => n496, D => n3002, Z => 
                           n3692);
   U3677 : NR4 port map( A => n3696, B => n3697, C => n3698, D => n3699, Z => 
                           n3685);
   U3678 : AO4 port map( A => n1568, B => n3007, C => n497, D => n3008, Z => 
                           n3699);
   U3679 : AO4 port map( A => n1569, B => n3009, C => n498, D => n3010, Z => 
                           n3698);
   U3680 : AO4 port map( A => n1570, B => n3011, C => n499, D => n3012, Z => 
                           n3697);
   U3681 : AO4 port map( A => n1571, B => n3013, C => n500, D => n3014, Z => 
                           n3696);
   U3682 : NR4 port map( A => n3700, B => n3701, C => n3702, D => n3703, Z => 
                           n3684);
   U3683 : AO4 port map( A => n1572, B => n3019, C => n501, D => n3020, Z => 
                           n3703);
   U3684 : AO4 port map( A => n1573, B => n3021, C => n502, D => n3022, Z => 
                           n3702);
   U3685 : AO4 port map( A => n1574, B => n3023, C => n503, D => n3024, Z => 
                           n3701);
   U3686 : AO4 port map( A => n1575, B => n3025, C => n504, D => n3026, Z => 
                           n3700);
   U3687 : ND4 port map( A => n3704, B => n3705, C => n3706, D => n3707, Z => 
                           n3682);
   U3688 : NR4 port map( A => n3708, B => n3709, C => n3710, D => n3711, Z => 
                           n3707);
   U3689 : AO4 port map( A => n1576, B => n3035, C => n505, D => n3036, Z => 
                           n3711);
   U3690 : AO4 port map( A => n1577, B => n3037, C => n506, D => n3038, Z => 
                           n3710);
   U3691 : AO4 port map( A => n1578, B => n3039, C => n507, D => n3040, Z => 
                           n3709);
   U3692 : AO4 port map( A => n1579, B => n3041, C => n508, D => n3042, Z => 
                           n3708);
   U3693 : NR4 port map( A => n3712, B => n3713, C => n3714, D => n3715, Z => 
                           n3706);
   U3694 : AO4 port map( A => n1580, B => n3047, C => n509, D => n3048, Z => 
                           n3715);
   U3695 : AO4 port map( A => n1581, B => n3049, C => n510, D => n3050, Z => 
                           n3714);
   U3696 : AO4 port map( A => n1582, B => n3051, C => n511, D => n3052, Z => 
                           n3713);
   U3697 : AO4 port map( A => n1583, B => n3053, C => n512, D => n3054, Z => 
                           n3712);
   U3698 : NR4 port map( A => n3716, B => n3717, C => n3718, D => n3719, Z => 
                           n3705);
   U3699 : AO4 port map( A => n1584, B => n3059, C => n513, D => n3060, Z => 
                           n3719);
   U3700 : AO4 port map( A => n1585, B => n3061, C => n514, D => n3062, Z => 
                           n3718);
   U3701 : AO4 port map( A => n1586, B => n3063, C => n515, D => n3064, Z => 
                           n3717);
   U3702 : AO4 port map( A => n1587, B => n3065, C => n516, D => n3066, Z => 
                           n3716);
   U3703 : NR4 port map( A => n3720, B => n3721, C => n3722, D => n3723, Z => 
                           n3704);
   U3704 : AO4 port map( A => n1588, B => n3071, C => n517, D => n3072, Z => 
                           n3723);
   U3705 : AO4 port map( A => n1589, B => n3073, C => n518, D => n3074, Z => 
                           n3722);
   U3706 : AO4 port map( A => n1590, B => n3075, C => n519, D => n3076, Z => 
                           n3721);
   U3707 : AO4 port map( A => n1591, B => n3077, C => n520, D => n3078, Z => 
                           n3720);
   U3708 : MUX21L port map( A => n1049, B => n3724, S => CE_I, Z => n4564);
   U3709 : NR2 port map( A => n3725, B => n3726, Z => n3724);
   U3710 : ND4 port map( A => n3727, B => n3728, C => n3729, D => n3730, Z => 
                           n3726);
   U3711 : NR4 port map( A => n3731, B => n3732, C => n3733, D => n3734, Z => 
                           n3730);
   U3712 : AO4 port map( A => n1592, B => n2983, C => n521, D => n2984, Z => 
                           n3734);
   U3713 : AO4 port map( A => n1593, B => n2985, C => n522, D => n2986, Z => 
                           n3733);
   U3714 : AO4 port map( A => n1594, B => n2987, C => n523, D => n2988, Z => 
                           n3732);
   U3715 : AO4 port map( A => n1595, B => n2989, C => n524, D => n2990, Z => 
                           n3731);
   U3716 : NR4 port map( A => n3735, B => n3736, C => n3737, D => n3738, Z => 
                           n3729);
   U3717 : AO4 port map( A => n1596, B => n2995, C => n525, D => n2996, Z => 
                           n3738);
   U3718 : AO4 port map( A => n1597, B => n2997, C => n526, D => n2998, Z => 
                           n3737);
   U3719 : AO4 port map( A => n1598, B => n2999, C => n527, D => n3000, Z => 
                           n3736);
   U3720 : AO4 port map( A => n1599, B => n3001, C => n528, D => n3002, Z => 
                           n3735);
   U3721 : NR4 port map( A => n3739, B => n3740, C => n3741, D => n3742, Z => 
                           n3728);
   U3722 : AO4 port map( A => n1600, B => n3007, C => n529, D => n3008, Z => 
                           n3742);
   U3723 : AO4 port map( A => n1601, B => n3009, C => n530, D => n3010, Z => 
                           n3741);
   U3724 : AO4 port map( A => n1602, B => n3011, C => n531, D => n3012, Z => 
                           n3740);
   U3725 : AO4 port map( A => n1603, B => n3013, C => n532, D => n3014, Z => 
                           n3739);
   U3726 : NR4 port map( A => n3743, B => n3744, C => n3745, D => n3746, Z => 
                           n3727);
   U3727 : AO4 port map( A => n1604, B => n3019, C => n533, D => n3020, Z => 
                           n3746);
   U3728 : AO4 port map( A => n1605, B => n3021, C => n534, D => n3022, Z => 
                           n3745);
   U3729 : AO4 port map( A => n1606, B => n3023, C => n535, D => n3024, Z => 
                           n3744);
   U3730 : AO4 port map( A => n1607, B => n3025, C => n536, D => n3026, Z => 
                           n3743);
   U3731 : ND4 port map( A => n3747, B => n3748, C => n3749, D => n3750, Z => 
                           n3725);
   U3732 : NR4 port map( A => n3751, B => n3752, C => n3753, D => n3754, Z => 
                           n3750);
   U3733 : AO4 port map( A => n1608, B => n3035, C => n537, D => n3036, Z => 
                           n3754);
   U3734 : AO4 port map( A => n1609, B => n3037, C => n538, D => n3038, Z => 
                           n3753);
   U3735 : AO4 port map( A => n1610, B => n3039, C => n539, D => n3040, Z => 
                           n3752);
   U3736 : AO4 port map( A => n1611, B => n3041, C => n540, D => n3042, Z => 
                           n3751);
   U3737 : NR4 port map( A => n3755, B => n3756, C => n3757, D => n3758, Z => 
                           n3749);
   U3738 : AO4 port map( A => n1612, B => n3047, C => n541, D => n3048, Z => 
                           n3758);
   U3739 : AO4 port map( A => n1613, B => n3049, C => n542, D => n3050, Z => 
                           n3757);
   U3740 : AO4 port map( A => n1614, B => n3051, C => n543, D => n3052, Z => 
                           n3756);
   U3741 : AO4 port map( A => n1615, B => n3053, C => n544, D => n3054, Z => 
                           n3755);
   U3742 : NR4 port map( A => n3759, B => n3760, C => n3761, D => n3762, Z => 
                           n3748);
   U3743 : AO4 port map( A => n1616, B => n3059, C => n545, D => n3060, Z => 
                           n3762);
   U3744 : AO4 port map( A => n1617, B => n3061, C => n546, D => n3062, Z => 
                           n3761);
   U3745 : AO4 port map( A => n1618, B => n3063, C => n547, D => n3064, Z => 
                           n3760);
   U3746 : AO4 port map( A => n1619, B => n3065, C => n548, D => n3066, Z => 
                           n3759);
   U3747 : NR4 port map( A => n3763, B => n3764, C => n3765, D => n3766, Z => 
                           n3747);
   U3748 : AO4 port map( A => n1620, B => n3071, C => n549, D => n3072, Z => 
                           n3766);
   U3749 : AO4 port map( A => n1621, B => n3073, C => n550, D => n3074, Z => 
                           n3765);
   U3750 : AO4 port map( A => n1622, B => n3075, C => n551, D => n3076, Z => 
                           n3764);
   U3751 : AO4 port map( A => n1623, B => n3077, C => n552, D => n3078, Z => 
                           n3763);
   U3752 : MUX21L port map( A => n1055, B => n3767, S => CE_I, Z => n4563);
   U3753 : NR2 port map( A => n3768, B => n3769, Z => n3767);
   U3754 : ND4 port map( A => n3770, B => n3771, C => n3772, D => n3773, Z => 
                           n3769);
   U3755 : NR4 port map( A => n3774, B => n3775, C => n3776, D => n3777, Z => 
                           n3773);
   U3756 : AO4 port map( A => n1624, B => n2983, C => n553, D => n2984, Z => 
                           n3777);
   U3757 : AO4 port map( A => n1625, B => n2985, C => n554, D => n2986, Z => 
                           n3776);
   U3758 : AO4 port map( A => n1626, B => n2987, C => n555, D => n2988, Z => 
                           n3775);
   U3759 : AO4 port map( A => n1627, B => n2989, C => n556, D => n2990, Z => 
                           n3774);
   U3760 : NR4 port map( A => n3778, B => n3779, C => n3780, D => n3781, Z => 
                           n3772);
   U3761 : AO4 port map( A => n1628, B => n2995, C => n557, D => n2996, Z => 
                           n3781);
   U3762 : AO4 port map( A => n1629, B => n2997, C => n558, D => n2998, Z => 
                           n3780);
   U3763 : AO4 port map( A => n1630, B => n2999, C => n559, D => n3000, Z => 
                           n3779);
   U3764 : AO4 port map( A => n1631, B => n3001, C => n560, D => n3002, Z => 
                           n3778);
   U3765 : NR4 port map( A => n3782, B => n3783, C => n3784, D => n3785, Z => 
                           n3771);
   U3766 : AO4 port map( A => n1632, B => n3007, C => n561, D => n3008, Z => 
                           n3785);
   U3767 : AO4 port map( A => n1633, B => n3009, C => n562, D => n3010, Z => 
                           n3784);
   U3768 : AO4 port map( A => n1634, B => n3011, C => n563, D => n3012, Z => 
                           n3783);
   U3769 : AO4 port map( A => n1635, B => n3013, C => n564, D => n3014, Z => 
                           n3782);
   U3770 : NR4 port map( A => n3786, B => n3787, C => n3788, D => n3789, Z => 
                           n3770);
   U3771 : AO4 port map( A => n1636, B => n3019, C => n565, D => n3020, Z => 
                           n3789);
   U3772 : AO4 port map( A => n1637, B => n3021, C => n566, D => n3022, Z => 
                           n3788);
   U3773 : AO4 port map( A => n1638, B => n3023, C => n567, D => n3024, Z => 
                           n3787);
   U3774 : AO4 port map( A => n1639, B => n3025, C => n568, D => n3026, Z => 
                           n3786);
   U3775 : ND4 port map( A => n3790, B => n3791, C => n3792, D => n3793, Z => 
                           n3768);
   U3776 : NR4 port map( A => n3794, B => n3795, C => n3796, D => n3797, Z => 
                           n3793);
   U3777 : AO4 port map( A => n1640, B => n3035, C => n569, D => n3036, Z => 
                           n3797);
   U3778 : AO4 port map( A => n1641, B => n3037, C => n570, D => n3038, Z => 
                           n3796);
   U3779 : AO4 port map( A => n1642, B => n3039, C => n571, D => n3040, Z => 
                           n3795);
   U3780 : AO4 port map( A => n1643, B => n3041, C => n572, D => n3042, Z => 
                           n3794);
   U3781 : NR4 port map( A => n3798, B => n3799, C => n3800, D => n3801, Z => 
                           n3792);
   U3782 : AO4 port map( A => n1644, B => n3047, C => n573, D => n3048, Z => 
                           n3801);
   U3783 : AO4 port map( A => n1645, B => n3049, C => n574, D => n3050, Z => 
                           n3800);
   U3784 : AO4 port map( A => n1646, B => n3051, C => n575, D => n3052, Z => 
                           n3799);
   U3785 : AO4 port map( A => n1647, B => n3053, C => n576, D => n3054, Z => 
                           n3798);
   U3786 : NR4 port map( A => n3802, B => n3803, C => n3804, D => n3805, Z => 
                           n3791);
   U3787 : AO4 port map( A => n1648, B => n3059, C => n577, D => n3060, Z => 
                           n3805);
   U3788 : AO4 port map( A => n1649, B => n3061, C => n578, D => n3062, Z => 
                           n3804);
   U3789 : AO4 port map( A => n1650, B => n3063, C => n579, D => n3064, Z => 
                           n3803);
   U3790 : AO4 port map( A => n1651, B => n3065, C => n580, D => n3066, Z => 
                           n3802);
   U3791 : NR4 port map( A => n3806, B => n3807, C => n3808, D => n3809, Z => 
                           n3790);
   U3792 : AO4 port map( A => n1652, B => n3071, C => n581, D => n3072, Z => 
                           n3809);
   U3793 : AO4 port map( A => n1653, B => n3073, C => n582, D => n3074, Z => 
                           n3808);
   U3794 : AO4 port map( A => n1654, B => n3075, C => n583, D => n3076, Z => 
                           n3807);
   U3795 : AO4 port map( A => n1655, B => n3077, C => n584, D => n3078, Z => 
                           n3806);
   U3796 : MUX21L port map( A => n1064, B => n3810, S => CE_I, Z => n4562);
   U3797 : NR2 port map( A => n3811, B => n3812, Z => n3810);
   U3798 : ND4 port map( A => n3813, B => n3814, C => n3815, D => n3816, Z => 
                           n3812);
   U3799 : NR4 port map( A => n3817, B => n3818, C => n3819, D => n3820, Z => 
                           n3816);
   U3800 : AO4 port map( A => n1656, B => n2983, C => n585, D => n2984, Z => 
                           n3820);
   U3801 : AO4 port map( A => n1657, B => n2985, C => n586, D => n2986, Z => 
                           n3819);
   U3802 : AO4 port map( A => n1658, B => n2987, C => n587, D => n2988, Z => 
                           n3818);
   U3803 : AO4 port map( A => n1659, B => n2989, C => n588, D => n2990, Z => 
                           n3817);
   U3804 : NR4 port map( A => n3821, B => n3822, C => n3823, D => n3824, Z => 
                           n3815);
   U3805 : AO4 port map( A => n1660, B => n2995, C => n589, D => n2996, Z => 
                           n3824);
   U3806 : AO4 port map( A => n1661, B => n2997, C => n590, D => n2998, Z => 
                           n3823);
   U3807 : AO4 port map( A => n1662, B => n2999, C => n591, D => n3000, Z => 
                           n3822);
   U3808 : AO4 port map( A => n1663, B => n3001, C => n592, D => n3002, Z => 
                           n3821);
   U3809 : NR4 port map( A => n3825, B => n3826, C => n3827, D => n3828, Z => 
                           n3814);
   U3810 : AO4 port map( A => n1664, B => n3007, C => n593, D => n3008, Z => 
                           n3828);
   U3811 : AO4 port map( A => n1665, B => n3009, C => n594, D => n3010, Z => 
                           n3827);
   U3812 : AO4 port map( A => n1666, B => n3011, C => n595, D => n3012, Z => 
                           n3826);
   U3813 : AO4 port map( A => n1667, B => n3013, C => n596, D => n3014, Z => 
                           n3825);
   U3814 : NR4 port map( A => n3829, B => n3830, C => n3831, D => n3832, Z => 
                           n3813);
   U3815 : AO4 port map( A => n1668, B => n3019, C => n597, D => n3020, Z => 
                           n3832);
   U3816 : AO4 port map( A => n1669, B => n3021, C => n598, D => n3022, Z => 
                           n3831);
   U3817 : AO4 port map( A => n1670, B => n3023, C => n599, D => n3024, Z => 
                           n3830);
   U3818 : AO4 port map( A => n1671, B => n3025, C => n600, D => n3026, Z => 
                           n3829);
   U3819 : ND4 port map( A => n3833, B => n3834, C => n3835, D => n3836, Z => 
                           n3811);
   U3820 : NR4 port map( A => n3837, B => n3838, C => n3839, D => n3840, Z => 
                           n3836);
   U3821 : AO4 port map( A => n1672, B => n3035, C => n601, D => n3036, Z => 
                           n3840);
   U3822 : AO4 port map( A => n1673, B => n3037, C => n602, D => n3038, Z => 
                           n3839);
   U3823 : AO4 port map( A => n1674, B => n3039, C => n603, D => n3040, Z => 
                           n3838);
   U3824 : AO4 port map( A => n1675, B => n3041, C => n604, D => n3042, Z => 
                           n3837);
   U3825 : NR4 port map( A => n3841, B => n3842, C => n3843, D => n3844, Z => 
                           n3835);
   U3826 : AO4 port map( A => n1676, B => n3047, C => n605, D => n3048, Z => 
                           n3844);
   U3827 : AO4 port map( A => n1677, B => n3049, C => n606, D => n3050, Z => 
                           n3843);
   U3828 : AO4 port map( A => n1678, B => n3051, C => n607, D => n3052, Z => 
                           n3842);
   U3829 : AO4 port map( A => n1679, B => n3053, C => n608, D => n3054, Z => 
                           n3841);
   U3830 : NR4 port map( A => n3845, B => n3846, C => n3847, D => n3848, Z => 
                           n3834);
   U3831 : AO4 port map( A => n1680, B => n3059, C => n609, D => n3060, Z => 
                           n3848);
   U3832 : AO4 port map( A => n1681, B => n3061, C => n610, D => n3062, Z => 
                           n3847);
   U3833 : AO4 port map( A => n1682, B => n3063, C => n611, D => n3064, Z => 
                           n3846);
   U3834 : AO4 port map( A => n1683, B => n3065, C => n612, D => n3066, Z => 
                           n3845);
   U3835 : NR4 port map( A => n3849, B => n3850, C => n3851, D => n3852, Z => 
                           n3833);
   U3836 : AO4 port map( A => n1684, B => n3071, C => n613, D => n3072, Z => 
                           n3852);
   U3837 : AO4 port map( A => n1685, B => n3073, C => n614, D => n3074, Z => 
                           n3851);
   U3838 : AO4 port map( A => n1686, B => n3075, C => n615, D => n3076, Z => 
                           n3850);
   U3839 : AO4 port map( A => n1687, B => n3077, C => n616, D => n3078, Z => 
                           n3849);
   U3840 : MUX21L port map( A => n1072, B => n3853, S => CE_I, Z => n4561);
   U3841 : NR2 port map( A => n3854, B => n3855, Z => n3853);
   U3842 : ND4 port map( A => n3856, B => n3857, C => n3858, D => n3859, Z => 
                           n3855);
   U3843 : NR4 port map( A => n3860, B => n3861, C => n3862, D => n3863, Z => 
                           n3859);
   U3844 : AO4 port map( A => n1688, B => n2983, C => n617, D => n2984, Z => 
                           n3863);
   U3845 : AO4 port map( A => n1689, B => n2985, C => n618, D => n2986, Z => 
                           n3862);
   U3846 : AO4 port map( A => n1690, B => n2987, C => n619, D => n2988, Z => 
                           n3861);
   U3847 : AO4 port map( A => n1691, B => n2989, C => n620, D => n2990, Z => 
                           n3860);
   U3848 : NR4 port map( A => n3864, B => n3865, C => n3866, D => n3867, Z => 
                           n3858);
   U3849 : AO4 port map( A => n1692, B => n2995, C => n621, D => n2996, Z => 
                           n3867);
   U3850 : AO4 port map( A => n1693, B => n2997, C => n622, D => n2998, Z => 
                           n3866);
   U3851 : AO4 port map( A => n1694, B => n2999, C => n623, D => n3000, Z => 
                           n3865);
   U3852 : AO4 port map( A => n1695, B => n3001, C => n624, D => n3002, Z => 
                           n3864);
   U3853 : NR4 port map( A => n3868, B => n3869, C => n3870, D => n3871, Z => 
                           n3857);
   U3854 : AO4 port map( A => n1696, B => n3007, C => n625, D => n3008, Z => 
                           n3871);
   U3855 : AO4 port map( A => n1697, B => n3009, C => n626, D => n3010, Z => 
                           n3870);
   U3856 : AO4 port map( A => n1698, B => n3011, C => n627, D => n3012, Z => 
                           n3869);
   U3857 : AO4 port map( A => n1699, B => n3013, C => n628, D => n3014, Z => 
                           n3868);
   U3858 : NR4 port map( A => n3872, B => n3873, C => n3874, D => n3875, Z => 
                           n3856);
   U3859 : AO4 port map( A => n1700, B => n3019, C => n629, D => n3020, Z => 
                           n3875);
   U3860 : AO4 port map( A => n1701, B => n3021, C => n630, D => n3022, Z => 
                           n3874);
   U3861 : AO4 port map( A => n1702, B => n3023, C => n631, D => n3024, Z => 
                           n3873);
   U3862 : AO4 port map( A => n1703, B => n3025, C => n632, D => n3026, Z => 
                           n3872);
   U3863 : ND4 port map( A => n3876, B => n3877, C => n3878, D => n3879, Z => 
                           n3854);
   U3864 : NR4 port map( A => n3880, B => n3881, C => n3882, D => n3883, Z => 
                           n3879);
   U3865 : AO4 port map( A => n1704, B => n3035, C => n633, D => n3036, Z => 
                           n3883);
   U3866 : AO4 port map( A => n1705, B => n3037, C => n634, D => n3038, Z => 
                           n3882);
   U3867 : AO4 port map( A => n1706, B => n3039, C => n635, D => n3040, Z => 
                           n3881);
   U3868 : AO4 port map( A => n1707, B => n3041, C => n636, D => n3042, Z => 
                           n3880);
   U3869 : NR4 port map( A => n3884, B => n3885, C => n3886, D => n3887, Z => 
                           n3878);
   U3870 : AO4 port map( A => n1708, B => n3047, C => n637, D => n3048, Z => 
                           n3887);
   U3871 : AO4 port map( A => n1709, B => n3049, C => n638, D => n3050, Z => 
                           n3886);
   U3872 : AO4 port map( A => n1710, B => n3051, C => n639, D => n3052, Z => 
                           n3885);
   U3873 : AO4 port map( A => n1711, B => n3053, C => n640, D => n3054, Z => 
                           n3884);
   U3874 : NR4 port map( A => n3888, B => n3889, C => n3890, D => n3891, Z => 
                           n3877);
   U3875 : AO4 port map( A => n1712, B => n3059, C => n641, D => n3060, Z => 
                           n3891);
   U3876 : AO4 port map( A => n1713, B => n3061, C => n642, D => n3062, Z => 
                           n3890);
   U3877 : AO4 port map( A => n1714, B => n3063, C => n643, D => n3064, Z => 
                           n3889);
   U3878 : AO4 port map( A => n1715, B => n3065, C => n644, D => n3066, Z => 
                           n3888);
   U3879 : NR4 port map( A => n3892, B => n3893, C => n3894, D => n3895, Z => 
                           n3876);
   U3880 : AO4 port map( A => n1716, B => n3071, C => n645, D => n3072, Z => 
                           n3895);
   U3881 : AO4 port map( A => n1717, B => n3073, C => n646, D => n3074, Z => 
                           n3894);
   U3882 : AO4 port map( A => n1718, B => n3075, C => n647, D => n3076, Z => 
                           n3893);
   U3883 : AO4 port map( A => n1719, B => n3077, C => n648, D => n3078, Z => 
                           n3892);
   U3884 : MUX21L port map( A => n1052, B => n3896, S => CE_I, Z => n4560);
   U3885 : NR2 port map( A => n3897, B => n3898, Z => n3896);
   U3886 : ND4 port map( A => n3899, B => n3900, C => n3901, D => n3902, Z => 
                           n3898);
   U3887 : NR4 port map( A => n3903, B => n3904, C => n3905, D => n3906, Z => 
                           n3902);
   U3888 : AO4 port map( A => n1720, B => n2983, C => n649, D => n2984, Z => 
                           n3906);
   U3889 : AO4 port map( A => n1721, B => n2985, C => n650, D => n2986, Z => 
                           n3905);
   U3890 : AO4 port map( A => n1722, B => n2987, C => n651, D => n2988, Z => 
                           n3904);
   U3891 : AO4 port map( A => n1723, B => n2989, C => n652, D => n2990, Z => 
                           n3903);
   U3892 : NR4 port map( A => n3907, B => n3908, C => n3909, D => n3910, Z => 
                           n3901);
   U3893 : AO4 port map( A => n1724, B => n2995, C => n653, D => n2996, Z => 
                           n3910);
   U3894 : AO4 port map( A => n1725, B => n2997, C => n654, D => n2998, Z => 
                           n3909);
   U3895 : AO4 port map( A => n1726, B => n2999, C => n655, D => n3000, Z => 
                           n3908);
   U3896 : AO4 port map( A => n1727, B => n3001, C => n656, D => n3002, Z => 
                           n3907);
   U3897 : NR4 port map( A => n3911, B => n3912, C => n3913, D => n3914, Z => 
                           n3900);
   U3898 : AO4 port map( A => n1728, B => n3007, C => n657, D => n3008, Z => 
                           n3914);
   U3899 : AO4 port map( A => n1729, B => n3009, C => n658, D => n3010, Z => 
                           n3913);
   U3900 : AO4 port map( A => n1730, B => n3011, C => n659, D => n3012, Z => 
                           n3912);
   U3901 : AO4 port map( A => n1731, B => n3013, C => n660, D => n3014, Z => 
                           n3911);
   U3902 : NR4 port map( A => n3915, B => n3916, C => n3917, D => n3918, Z => 
                           n3899);
   U3903 : AO4 port map( A => n1732, B => n3019, C => n661, D => n3020, Z => 
                           n3918);
   U3904 : AO4 port map( A => n1733, B => n3021, C => n662, D => n3022, Z => 
                           n3917);
   U3905 : AO4 port map( A => n1734, B => n3023, C => n663, D => n3024, Z => 
                           n3916);
   U3906 : AO4 port map( A => n1735, B => n3025, C => n664, D => n3026, Z => 
                           n3915);
   U3907 : ND4 port map( A => n3919, B => n3920, C => n3921, D => n3922, Z => 
                           n3897);
   U3908 : NR4 port map( A => n3923, B => n3924, C => n3925, D => n3926, Z => 
                           n3922);
   U3909 : AO4 port map( A => n1736, B => n3035, C => n665, D => n3036, Z => 
                           n3926);
   U3910 : AO4 port map( A => n1737, B => n3037, C => n666, D => n3038, Z => 
                           n3925);
   U3911 : AO4 port map( A => n1738, B => n3039, C => n667, D => n3040, Z => 
                           n3924);
   U3912 : AO4 port map( A => n1739, B => n3041, C => n668, D => n3042, Z => 
                           n3923);
   U3913 : NR4 port map( A => n3927, B => n3928, C => n3929, D => n3930, Z => 
                           n3921);
   U3914 : AO4 port map( A => n1740, B => n3047, C => n669, D => n3048, Z => 
                           n3930);
   U3915 : AO4 port map( A => n1741, B => n3049, C => n670, D => n3050, Z => 
                           n3929);
   U3916 : AO4 port map( A => n1742, B => n3051, C => n671, D => n3052, Z => 
                           n3928);
   U3917 : AO4 port map( A => n1743, B => n3053, C => n672, D => n3054, Z => 
                           n3927);
   U3918 : NR4 port map( A => n3931, B => n3932, C => n3933, D => n3934, Z => 
                           n3920);
   U3919 : AO4 port map( A => n1744, B => n3059, C => n673, D => n3060, Z => 
                           n3934);
   U3920 : AO4 port map( A => n1745, B => n3061, C => n674, D => n3062, Z => 
                           n3933);
   U3921 : AO4 port map( A => n1746, B => n3063, C => n675, D => n3064, Z => 
                           n3932);
   U3922 : AO4 port map( A => n1747, B => n3065, C => n676, D => n3066, Z => 
                           n3931);
   U3923 : NR4 port map( A => n3935, B => n3936, C => n3937, D => n3938, Z => 
                           n3919);
   U3924 : AO4 port map( A => n1748, B => n3071, C => n677, D => n3072, Z => 
                           n3938);
   U3925 : AO4 port map( A => n1749, B => n3073, C => n678, D => n3074, Z => 
                           n3937);
   U3926 : AO4 port map( A => n1750, B => n3075, C => n679, D => n3076, Z => 
                           n3936);
   U3927 : AO4 port map( A => n1751, B => n3077, C => n680, D => n3078, Z => 
                           n3935);
   U3928 : MUX21L port map( A => n1056, B => n3939, S => CE_I, Z => n4559);
   U3929 : NR2 port map( A => n3940, B => n3941, Z => n3939);
   U3930 : ND4 port map( A => n3942, B => n3943, C => n3944, D => n3945, Z => 
                           n3941);
   U3931 : NR4 port map( A => n3946, B => n3947, C => n3948, D => n3949, Z => 
                           n3945);
   U3932 : AO4 port map( A => n1752, B => n2983, C => n681, D => n2984, Z => 
                           n3949);
   U3933 : AO4 port map( A => n1753, B => n2985, C => n682, D => n2986, Z => 
                           n3948);
   U3934 : AO4 port map( A => n1754, B => n2987, C => n683, D => n2988, Z => 
                           n3947);
   U3935 : AO4 port map( A => n1755, B => n2989, C => n684, D => n2990, Z => 
                           n3946);
   U3936 : NR4 port map( A => n3950, B => n3951, C => n3952, D => n3953, Z => 
                           n3944);
   U3937 : AO4 port map( A => n1756, B => n2995, C => n685, D => n2996, Z => 
                           n3953);
   U3938 : AO4 port map( A => n1757, B => n2997, C => n686, D => n2998, Z => 
                           n3952);
   U3939 : AO4 port map( A => n1758, B => n2999, C => n687, D => n3000, Z => 
                           n3951);
   U3940 : AO4 port map( A => n1759, B => n3001, C => n688, D => n3002, Z => 
                           n3950);
   U3941 : NR4 port map( A => n3954, B => n3955, C => n3956, D => n3957, Z => 
                           n3943);
   U3942 : AO4 port map( A => n1760, B => n3007, C => n689, D => n3008, Z => 
                           n3957);
   U3943 : AO4 port map( A => n1761, B => n3009, C => n690, D => n3010, Z => 
                           n3956);
   U3944 : AO4 port map( A => n1762, B => n3011, C => n691, D => n3012, Z => 
                           n3955);
   U3945 : AO4 port map( A => n1763, B => n3013, C => n692, D => n3014, Z => 
                           n3954);
   U3946 : NR4 port map( A => n3958, B => n3959, C => n3960, D => n3961, Z => 
                           n3942);
   U3947 : AO4 port map( A => n1764, B => n3019, C => n693, D => n3020, Z => 
                           n3961);
   U3948 : AO4 port map( A => n1765, B => n3021, C => n694, D => n3022, Z => 
                           n3960);
   U3949 : AO4 port map( A => n1766, B => n3023, C => n695, D => n3024, Z => 
                           n3959);
   U3950 : AO4 port map( A => n1767, B => n3025, C => n696, D => n3026, Z => 
                           n3958);
   U3951 : ND4 port map( A => n3962, B => n3963, C => n3964, D => n3965, Z => 
                           n3940);
   U3952 : NR4 port map( A => n3966, B => n3967, C => n3968, D => n3969, Z => 
                           n3965);
   U3953 : AO4 port map( A => n1768, B => n3035, C => n697, D => n3036, Z => 
                           n3969);
   U3954 : AO4 port map( A => n1769, B => n3037, C => n698, D => n3038, Z => 
                           n3968);
   U3955 : AO4 port map( A => n1770, B => n3039, C => n699, D => n3040, Z => 
                           n3967);
   U3956 : AO4 port map( A => n1771, B => n3041, C => n700, D => n3042, Z => 
                           n3966);
   U3957 : NR4 port map( A => n3970, B => n3971, C => n3972, D => n3973, Z => 
                           n3964);
   U3958 : AO4 port map( A => n1772, B => n3047, C => n701, D => n3048, Z => 
                           n3973);
   U3959 : AO4 port map( A => n1773, B => n3049, C => n702, D => n3050, Z => 
                           n3972);
   U3960 : AO4 port map( A => n1774, B => n3051, C => n703, D => n3052, Z => 
                           n3971);
   U3961 : AO4 port map( A => n1775, B => n3053, C => n704, D => n3054, Z => 
                           n3970);
   U3962 : NR4 port map( A => n3974, B => n3975, C => n3976, D => n3977, Z => 
                           n3963);
   U3963 : AO4 port map( A => n1776, B => n3059, C => n705, D => n3060, Z => 
                           n3977);
   U3964 : AO4 port map( A => n1777, B => n3061, C => n706, D => n3062, Z => 
                           n3976);
   U3965 : AO4 port map( A => n1778, B => n3063, C => n707, D => n3064, Z => 
                           n3975);
   U3966 : AO4 port map( A => n1779, B => n3065, C => n708, D => n3066, Z => 
                           n3974);
   U3967 : NR4 port map( A => n3978, B => n3979, C => n3980, D => n3981, Z => 
                           n3962);
   U3968 : AO4 port map( A => n1780, B => n3071, C => n709, D => n3072, Z => 
                           n3981);
   U3969 : AO4 port map( A => n1781, B => n3073, C => n710, D => n3074, Z => 
                           n3980);
   U3970 : AO4 port map( A => n1782, B => n3075, C => n711, D => n3076, Z => 
                           n3979);
   U3971 : AO4 port map( A => n1783, B => n3077, C => n712, D => n3078, Z => 
                           n3978);
   U3972 : MUX21L port map( A => n1065, B => n3982, S => CE_I, Z => n4558);
   U3973 : NR2 port map( A => n3983, B => n3984, Z => n3982);
   U3974 : ND4 port map( A => n3985, B => n3986, C => n3987, D => n3988, Z => 
                           n3984);
   U3975 : NR4 port map( A => n3989, B => n3990, C => n3991, D => n3992, Z => 
                           n3988);
   U3976 : AO4 port map( A => n1784, B => n2983, C => n713, D => n2984, Z => 
                           n3992);
   U3977 : AO4 port map( A => n1785, B => n2985, C => n714, D => n2986, Z => 
                           n3991);
   U3978 : AO4 port map( A => n1786, B => n2987, C => n715, D => n2988, Z => 
                           n3990);
   U3979 : AO4 port map( A => n1787, B => n2989, C => n716, D => n2990, Z => 
                           n3989);
   U3980 : NR4 port map( A => n3993, B => n3994, C => n3995, D => n3996, Z => 
                           n3987);
   U3981 : AO4 port map( A => n1788, B => n2995, C => n717, D => n2996, Z => 
                           n3996);
   U3982 : AO4 port map( A => n1789, B => n2997, C => n718, D => n2998, Z => 
                           n3995);
   U3983 : AO4 port map( A => n1790, B => n2999, C => n719, D => n3000, Z => 
                           n3994);
   U3984 : AO4 port map( A => n1791, B => n3001, C => n720, D => n3002, Z => 
                           n3993);
   U3985 : NR4 port map( A => n3997, B => n3998, C => n3999, D => n4000, Z => 
                           n3986);
   U3986 : AO4 port map( A => n1792, B => n3007, C => n721, D => n3008, Z => 
                           n4000);
   U3987 : AO4 port map( A => n1793, B => n3009, C => n722, D => n3010, Z => 
                           n3999);
   U3988 : AO4 port map( A => n1794, B => n3011, C => n723, D => n3012, Z => 
                           n3998);
   U3989 : AO4 port map( A => n1795, B => n3013, C => n724, D => n3014, Z => 
                           n3997);
   U3990 : NR4 port map( A => n4001, B => n4002, C => n4003, D => n4004, Z => 
                           n3985);
   U3991 : AO4 port map( A => n1796, B => n3019, C => n725, D => n3020, Z => 
                           n4004);
   U3992 : AO4 port map( A => n1797, B => n3021, C => n726, D => n3022, Z => 
                           n4003);
   U3993 : AO4 port map( A => n1798, B => n3023, C => n727, D => n3024, Z => 
                           n4002);
   U3994 : AO4 port map( A => n1799, B => n3025, C => n728, D => n3026, Z => 
                           n4001);
   U3995 : ND4 port map( A => n4005, B => n4006, C => n4007, D => n4008, Z => 
                           n3983);
   U3996 : NR4 port map( A => n4009, B => n4010, C => n4011, D => n4012, Z => 
                           n4008);
   U3997 : AO4 port map( A => n1800, B => n3035, C => n729, D => n3036, Z => 
                           n4012);
   U3998 : AO4 port map( A => n1801, B => n3037, C => n730, D => n3038, Z => 
                           n4011);
   U3999 : AO4 port map( A => n1802, B => n3039, C => n731, D => n3040, Z => 
                           n4010);
   U4000 : AO4 port map( A => n1803, B => n3041, C => n732, D => n3042, Z => 
                           n4009);
   U4001 : NR4 port map( A => n4013, B => n4014, C => n4015, D => n4016, Z => 
                           n4007);
   U4002 : AO4 port map( A => n1804, B => n3047, C => n733, D => n3048, Z => 
                           n4016);
   U4003 : AO4 port map( A => n1805, B => n3049, C => n734, D => n3050, Z => 
                           n4015);
   U4004 : AO4 port map( A => n1806, B => n3051, C => n735, D => n3052, Z => 
                           n4014);
   U4005 : AO4 port map( A => n1807, B => n3053, C => n736, D => n3054, Z => 
                           n4013);
   U4006 : NR4 port map( A => n4017, B => n4018, C => n4019, D => n4020, Z => 
                           n4006);
   U4007 : AO4 port map( A => n1808, B => n3059, C => n737, D => n3060, Z => 
                           n4020);
   U4008 : AO4 port map( A => n1809, B => n3061, C => n738, D => n3062, Z => 
                           n4019);
   U4009 : AO4 port map( A => n1810, B => n3063, C => n739, D => n3064, Z => 
                           n4018);
   U4010 : AO4 port map( A => n1811, B => n3065, C => n740, D => n3066, Z => 
                           n4017);
   U4011 : NR4 port map( A => n4021, B => n4022, C => n4023, D => n4024, Z => 
                           n4005);
   U4012 : AO4 port map( A => n1812, B => n3071, C => n741, D => n3072, Z => 
                           n4024);
   U4013 : AO4 port map( A => n1813, B => n3073, C => n742, D => n3074, Z => 
                           n4023);
   U4014 : AO4 port map( A => n1814, B => n3075, C => n743, D => n3076, Z => 
                           n4022);
   U4015 : AO4 port map( A => n1815, B => n3077, C => n744, D => n3078, Z => 
                           n4021);
   U4016 : MUX21L port map( A => n1073, B => n4025, S => CE_I, Z => n4557);
   U4017 : NR2 port map( A => n4026, B => n4027, Z => n4025);
   U4018 : ND4 port map( A => n4028, B => n4029, C => n4030, D => n4031, Z => 
                           n4027);
   U4019 : NR4 port map( A => n4032, B => n4033, C => n4034, D => n4035, Z => 
                           n4031);
   U4020 : AO4 port map( A => n1816, B => n2983, C => n745, D => n2984, Z => 
                           n4035);
   U4021 : AO4 port map( A => n1817, B => n2985, C => n746, D => n2986, Z => 
                           n4034);
   U4022 : AO4 port map( A => n1818, B => n2987, C => n747, D => n2988, Z => 
                           n4033);
   U4023 : AO4 port map( A => n1819, B => n2989, C => n748, D => n2990, Z => 
                           n4032);
   U4024 : NR4 port map( A => n4036, B => n4037, C => n4038, D => n4039, Z => 
                           n4030);
   U4025 : AO4 port map( A => n1820, B => n2995, C => n749, D => n2996, Z => 
                           n4039);
   U4026 : AO4 port map( A => n1821, B => n2997, C => n750, D => n2998, Z => 
                           n4038);
   U4027 : AO4 port map( A => n1822, B => n2999, C => n751, D => n3000, Z => 
                           n4037);
   U4028 : AO4 port map( A => n1823, B => n3001, C => n752, D => n3002, Z => 
                           n4036);
   U4029 : NR4 port map( A => n4040, B => n4041, C => n4042, D => n4043, Z => 
                           n4029);
   U4030 : AO4 port map( A => n1824, B => n3007, C => n753, D => n3008, Z => 
                           n4043);
   U4031 : AO4 port map( A => n1825, B => n3009, C => n754, D => n3010, Z => 
                           n4042);
   U4032 : AO4 port map( A => n1826, B => n3011, C => n755, D => n3012, Z => 
                           n4041);
   U4033 : AO4 port map( A => n1827, B => n3013, C => n756, D => n3014, Z => 
                           n4040);
   U4034 : NR4 port map( A => n4044, B => n4045, C => n4046, D => n4047, Z => 
                           n4028);
   U4035 : AO4 port map( A => n1828, B => n3019, C => n757, D => n3020, Z => 
                           n4047);
   U4036 : AO4 port map( A => n1829, B => n3021, C => n758, D => n3022, Z => 
                           n4046);
   U4037 : AO4 port map( A => n1830, B => n3023, C => n759, D => n3024, Z => 
                           n4045);
   U4038 : AO4 port map( A => n1831, B => n3025, C => n760, D => n3026, Z => 
                           n4044);
   U4039 : ND4 port map( A => n4048, B => n4049, C => n4050, D => n4051, Z => 
                           n4026);
   U4040 : NR4 port map( A => n4052, B => n4053, C => n4054, D => n4055, Z => 
                           n4051);
   U4041 : AO4 port map( A => n1832, B => n3035, C => n761, D => n3036, Z => 
                           n4055);
   U4042 : AO4 port map( A => n1833, B => n3037, C => n762, D => n3038, Z => 
                           n4054);
   U4043 : AO4 port map( A => n1834, B => n3039, C => n763, D => n3040, Z => 
                           n4053);
   U4044 : AO4 port map( A => n1835, B => n3041, C => n764, D => n3042, Z => 
                           n4052);
   U4045 : NR4 port map( A => n4056, B => n4057, C => n4058, D => n4059, Z => 
                           n4050);
   U4046 : AO4 port map( A => n1836, B => n3047, C => n765, D => n3048, Z => 
                           n4059);
   U4047 : AO4 port map( A => n1837, B => n3049, C => n766, D => n3050, Z => 
                           n4058);
   U4048 : AO4 port map( A => n1838, B => n3051, C => n767, D => n3052, Z => 
                           n4057);
   U4049 : AO4 port map( A => n1839, B => n3053, C => n768, D => n3054, Z => 
                           n4056);
   U4050 : NR4 port map( A => n4060, B => n4061, C => n4062, D => n4063, Z => 
                           n4049);
   U4051 : AO4 port map( A => n1840, B => n3059, C => n769, D => n3060, Z => 
                           n4063);
   U4052 : AO4 port map( A => n1841, B => n3061, C => n770, D => n3062, Z => 
                           n4062);
   U4053 : AO4 port map( A => n1842, B => n3063, C => n771, D => n3064, Z => 
                           n4061);
   U4054 : AO4 port map( A => n1843, B => n3065, C => n772, D => n3066, Z => 
                           n4060);
   U4055 : NR4 port map( A => n4064, B => n4065, C => n4066, D => n4067, Z => 
                           n4048);
   U4056 : AO4 port map( A => n1844, B => n3071, C => n773, D => n3072, Z => 
                           n4067);
   U4057 : AO4 port map( A => n1845, B => n3073, C => n774, D => n3074, Z => 
                           n4066);
   U4058 : AO4 port map( A => n1846, B => n3075, C => n775, D => n3076, Z => 
                           n4065);
   U4059 : AO4 port map( A => n1847, B => n3077, C => n776, D => n3078, Z => 
                           n4064);
   U4060 : MUX21L port map( A => n1063, B => n4068, S => CE_I, Z => n4556);
   U4061 : NR2 port map( A => n4069, B => n4070, Z => n4068);
   U4062 : ND4 port map( A => n4071, B => n4072, C => n4073, D => n4074, Z => 
                           n4070);
   U4063 : NR4 port map( A => n4075, B => n4076, C => n4077, D => n4078, Z => 
                           n4074);
   U4064 : AO4 port map( A => n1848, B => n2983, C => n777, D => n2984, Z => 
                           n4078);
   U4065 : AO4 port map( A => n1849, B => n2985, C => n778, D => n2986, Z => 
                           n4077);
   U4066 : AO4 port map( A => n1850, B => n2987, C => n779, D => n2988, Z => 
                           n4076);
   U4067 : AO4 port map( A => n1851, B => n2989, C => n780, D => n2990, Z => 
                           n4075);
   U4068 : NR4 port map( A => n4079, B => n4080, C => n4081, D => n4082, Z => 
                           n4073);
   U4069 : AO4 port map( A => n1852, B => n2995, C => n781, D => n2996, Z => 
                           n4082);
   U4070 : AO4 port map( A => n1853, B => n2997, C => n782, D => n2998, Z => 
                           n4081);
   U4071 : AO4 port map( A => n1854, B => n2999, C => n783, D => n3000, Z => 
                           n4080);
   U4072 : AO4 port map( A => n1855, B => n3001, C => n784, D => n3002, Z => 
                           n4079);
   U4073 : NR4 port map( A => n4083, B => n4084, C => n4085, D => n4086, Z => 
                           n4072);
   U4074 : AO4 port map( A => n1856, B => n3007, C => n785, D => n3008, Z => 
                           n4086);
   U4075 : AO4 port map( A => n1857, B => n3009, C => n786, D => n3010, Z => 
                           n4085);
   U4076 : AO4 port map( A => n1858, B => n3011, C => n787, D => n3012, Z => 
                           n4084);
   U4077 : AO4 port map( A => n1859, B => n3013, C => n788, D => n3014, Z => 
                           n4083);
   U4078 : NR4 port map( A => n4087, B => n4088, C => n4089, D => n4090, Z => 
                           n4071);
   U4079 : AO4 port map( A => n1860, B => n3019, C => n789, D => n3020, Z => 
                           n4090);
   U4080 : AO4 port map( A => n1861, B => n3021, C => n790, D => n3022, Z => 
                           n4089);
   U4081 : AO4 port map( A => n1862, B => n3023, C => n791, D => n3024, Z => 
                           n4088);
   U4082 : AO4 port map( A => n1863, B => n3025, C => n792, D => n3026, Z => 
                           n4087);
   U4083 : ND4 port map( A => n4091, B => n4092, C => n4093, D => n4094, Z => 
                           n4069);
   U4084 : NR4 port map( A => n4095, B => n4096, C => n4097, D => n4098, Z => 
                           n4094);
   U4085 : AO4 port map( A => n1864, B => n3035, C => n793, D => n3036, Z => 
                           n4098);
   U4086 : AO4 port map( A => n1865, B => n3037, C => n794, D => n3038, Z => 
                           n4097);
   U4087 : AO4 port map( A => n1866, B => n3039, C => n795, D => n3040, Z => 
                           n4096);
   U4088 : AO4 port map( A => n1867, B => n3041, C => n796, D => n3042, Z => 
                           n4095);
   U4089 : NR4 port map( A => n4099, B => n4100, C => n4101, D => n4102, Z => 
                           n4093);
   U4090 : AO4 port map( A => n1868, B => n3047, C => n797, D => n3048, Z => 
                           n4102);
   U4091 : AO4 port map( A => n1869, B => n3049, C => n798, D => n3050, Z => 
                           n4101);
   U4092 : AO4 port map( A => n1870, B => n3051, C => n799, D => n3052, Z => 
                           n4100);
   U4093 : AO4 port map( A => n1871, B => n3053, C => n800, D => n3054, Z => 
                           n4099);
   U4094 : NR4 port map( A => n4103, B => n4104, C => n4105, D => n4106, Z => 
                           n4092);
   U4095 : AO4 port map( A => n1872, B => n3059, C => n801, D => n3060, Z => 
                           n4106);
   U4096 : AO4 port map( A => n1873, B => n3061, C => n802, D => n3062, Z => 
                           n4105);
   U4097 : AO4 port map( A => n1874, B => n3063, C => n803, D => n3064, Z => 
                           n4104);
   U4098 : AO4 port map( A => n1875, B => n3065, C => n804, D => n3066, Z => 
                           n4103);
   U4099 : NR4 port map( A => n4107, B => n4108, C => n4109, D => n4110, Z => 
                           n4091);
   U4100 : AO4 port map( A => n1876, B => n3071, C => n805, D => n3072, Z => 
                           n4110);
   U4101 : AO4 port map( A => n1877, B => n3073, C => n806, D => n3074, Z => 
                           n4109);
   U4102 : AO4 port map( A => n1878, B => n3075, C => n807, D => n3076, Z => 
                           n4108);
   U4103 : AO4 port map( A => n1879, B => n3077, C => n808, D => n3078, Z => 
                           n4107);
   U4104 : MUX21L port map( A => n1057, B => n4111, S => CE_I, Z => n4555);
   U4105 : NR2 port map( A => n4112, B => n4113, Z => n4111);
   U4106 : ND4 port map( A => n4114, B => n4115, C => n4116, D => n4117, Z => 
                           n4113);
   U4107 : NR4 port map( A => n4118, B => n4119, C => n4120, D => n4121, Z => 
                           n4117);
   U4108 : AO4 port map( A => n1880, B => n2983, C => n809, D => n2984, Z => 
                           n4121);
   U4109 : AO4 port map( A => n1881, B => n2985, C => n810, D => n2986, Z => 
                           n4120);
   U4110 : AO4 port map( A => n1882, B => n2987, C => n811, D => n2988, Z => 
                           n4119);
   U4111 : AO4 port map( A => n1883, B => n2989, C => n812, D => n2990, Z => 
                           n4118);
   U4112 : NR4 port map( A => n4122, B => n4123, C => n4124, D => n4125, Z => 
                           n4116);
   U4113 : AO4 port map( A => n1884, B => n2995, C => n813, D => n2996, Z => 
                           n4125);
   U4114 : AO4 port map( A => n1885, B => n2997, C => n814, D => n2998, Z => 
                           n4124);
   U4115 : AO4 port map( A => n1886, B => n2999, C => n815, D => n3000, Z => 
                           n4123);
   U4116 : AO4 port map( A => n1887, B => n3001, C => n816, D => n3002, Z => 
                           n4122);
   U4117 : NR4 port map( A => n4126, B => n4127, C => n4128, D => n4129, Z => 
                           n4115);
   U4118 : AO4 port map( A => n1888, B => n3007, C => n817, D => n3008, Z => 
                           n4129);
   U4119 : AO4 port map( A => n1889, B => n3009, C => n818, D => n3010, Z => 
                           n4128);
   U4120 : AO4 port map( A => n1890, B => n3011, C => n819, D => n3012, Z => 
                           n4127);
   U4121 : AO4 port map( A => n1891, B => n3013, C => n820, D => n3014, Z => 
                           n4126);
   U4122 : NR4 port map( A => n4130, B => n4131, C => n4132, D => n4133, Z => 
                           n4114);
   U4123 : AO4 port map( A => n1892, B => n3019, C => n821, D => n3020, Z => 
                           n4133);
   U4124 : AO4 port map( A => n1893, B => n3021, C => n822, D => n3022, Z => 
                           n4132);
   U4125 : AO4 port map( A => n1894, B => n3023, C => n823, D => n3024, Z => 
                           n4131);
   U4126 : AO4 port map( A => n1895, B => n3025, C => n824, D => n3026, Z => 
                           n4130);
   U4127 : ND4 port map( A => n4134, B => n4135, C => n4136, D => n4137, Z => 
                           n4112);
   U4128 : NR4 port map( A => n4138, B => n4139, C => n4140, D => n4141, Z => 
                           n4137);
   U4129 : AO4 port map( A => n1896, B => n3035, C => n825, D => n3036, Z => 
                           n4141);
   U4130 : AO4 port map( A => n1897, B => n3037, C => n826, D => n3038, Z => 
                           n4140);
   U4131 : AO4 port map( A => n1898, B => n3039, C => n827, D => n3040, Z => 
                           n4139);
   U4132 : AO4 port map( A => n1899, B => n3041, C => n828, D => n3042, Z => 
                           n4138);
   U4133 : NR4 port map( A => n4142, B => n4143, C => n4144, D => n4145, Z => 
                           n4136);
   U4134 : AO4 port map( A => n1900, B => n3047, C => n829, D => n3048, Z => 
                           n4145);
   U4135 : AO4 port map( A => n1901, B => n3049, C => n830, D => n3050, Z => 
                           n4144);
   U4136 : AO4 port map( A => n1902, B => n3051, C => n831, D => n3052, Z => 
                           n4143);
   U4137 : AO4 port map( A => n1903, B => n3053, C => n832, D => n3054, Z => 
                           n4142);
   U4138 : NR4 port map( A => n4146, B => n4147, C => n4148, D => n4149, Z => 
                           n4135);
   U4139 : AO4 port map( A => n1904, B => n3059, C => n833, D => n3060, Z => 
                           n4149);
   U4140 : AO4 port map( A => n1905, B => n3061, C => n834, D => n3062, Z => 
                           n4148);
   U4141 : AO4 port map( A => n1906, B => n3063, C => n835, D => n3064, Z => 
                           n4147);
   U4142 : AO4 port map( A => n1907, B => n3065, C => n836, D => n3066, Z => 
                           n4146);
   U4143 : NR4 port map( A => n4150, B => n4151, C => n4152, D => n4153, Z => 
                           n4134);
   U4144 : AO4 port map( A => n1908, B => n3071, C => n837, D => n3072, Z => 
                           n4153);
   U4145 : AO4 port map( A => n1909, B => n3073, C => n838, D => n3074, Z => 
                           n4152);
   U4146 : AO4 port map( A => n1910, B => n3075, C => n839, D => n3076, Z => 
                           n4151);
   U4147 : AO4 port map( A => n1911, B => n3077, C => n840, D => n3078, Z => 
                           n4150);
   U4148 : MUX21L port map( A => n1066, B => n4154, S => CE_I, Z => n4554);
   U4149 : NR2 port map( A => n4155, B => n4156, Z => n4154);
   U4150 : ND4 port map( A => n4157, B => n4158, C => n4159, D => n4160, Z => 
                           n4156);
   U4151 : NR4 port map( A => n4161, B => n4162, C => n4163, D => n4164, Z => 
                           n4160);
   U4152 : AO4 port map( A => n1912, B => n2983, C => n841, D => n2984, Z => 
                           n4164);
   U4153 : AO4 port map( A => n1913, B => n2985, C => n842, D => n2986, Z => 
                           n4163);
   U4154 : AO4 port map( A => n1914, B => n2987, C => n843, D => n2988, Z => 
                           n4162);
   U4155 : AO4 port map( A => n1915, B => n2989, C => n844, D => n2990, Z => 
                           n4161);
   U4156 : NR4 port map( A => n4165, B => n4166, C => n4167, D => n4168, Z => 
                           n4159);
   U4157 : AO4 port map( A => n1916, B => n2995, C => n845, D => n2996, Z => 
                           n4168);
   U4158 : AO4 port map( A => n1917, B => n2997, C => n846, D => n2998, Z => 
                           n4167);
   U4159 : AO4 port map( A => n1918, B => n2999, C => n847, D => n3000, Z => 
                           n4166);
   U4160 : AO4 port map( A => n1919, B => n3001, C => n848, D => n3002, Z => 
                           n4165);
   U4161 : NR4 port map( A => n4169, B => n4170, C => n4171, D => n4172, Z => 
                           n4158);
   U4162 : AO4 port map( A => n1920, B => n3007, C => n849, D => n3008, Z => 
                           n4172);
   U4163 : AO4 port map( A => n1921, B => n3009, C => n850, D => n3010, Z => 
                           n4171);
   U4164 : AO4 port map( A => n1922, B => n3011, C => n851, D => n3012, Z => 
                           n4170);
   U4165 : AO4 port map( A => n1923, B => n3013, C => n852, D => n3014, Z => 
                           n4169);
   U4166 : NR4 port map( A => n4173, B => n4174, C => n4175, D => n4176, Z => 
                           n4157);
   U4167 : AO4 port map( A => n1924, B => n3019, C => n853, D => n3020, Z => 
                           n4176);
   U4168 : AO4 port map( A => n1925, B => n3021, C => n854, D => n3022, Z => 
                           n4175);
   U4169 : AO4 port map( A => n1926, B => n3023, C => n855, D => n3024, Z => 
                           n4174);
   U4170 : AO4 port map( A => n1927, B => n3025, C => n856, D => n3026, Z => 
                           n4173);
   U4171 : ND4 port map( A => n4177, B => n4178, C => n4179, D => n4180, Z => 
                           n4155);
   U4172 : NR4 port map( A => n4181, B => n4182, C => n4183, D => n4184, Z => 
                           n4180);
   U4173 : AO4 port map( A => n1928, B => n3035, C => n857, D => n3036, Z => 
                           n4184);
   U4174 : AO4 port map( A => n1929, B => n3037, C => n858, D => n3038, Z => 
                           n4183);
   U4175 : AO4 port map( A => n1930, B => n3039, C => n859, D => n3040, Z => 
                           n4182);
   U4176 : AO4 port map( A => n1931, B => n3041, C => n860, D => n3042, Z => 
                           n4181);
   U4177 : NR4 port map( A => n4185, B => n4186, C => n4187, D => n4188, Z => 
                           n4179);
   U4178 : AO4 port map( A => n1932, B => n3047, C => n861, D => n3048, Z => 
                           n4188);
   U4179 : AO4 port map( A => n1933, B => n3049, C => n862, D => n3050, Z => 
                           n4187);
   U4180 : AO4 port map( A => n1934, B => n3051, C => n863, D => n3052, Z => 
                           n4186);
   U4181 : AO4 port map( A => n1935, B => n3053, C => n864, D => n3054, Z => 
                           n4185);
   U4182 : NR4 port map( A => n4189, B => n4190, C => n4191, D => n4192, Z => 
                           n4178);
   U4183 : AO4 port map( A => n1936, B => n3059, C => n865, D => n3060, Z => 
                           n4192);
   U4184 : AO4 port map( A => n1937, B => n3061, C => n866, D => n3062, Z => 
                           n4191);
   U4185 : AO4 port map( A => n1938, B => n3063, C => n867, D => n3064, Z => 
                           n4190);
   U4186 : AO4 port map( A => n1939, B => n3065, C => n868, D => n3066, Z => 
                           n4189);
   U4187 : NR4 port map( A => n4193, B => n4194, C => n4195, D => n4196, Z => 
                           n4177);
   U4188 : AO4 port map( A => n1940, B => n3071, C => n869, D => n3072, Z => 
                           n4196);
   U4189 : AO4 port map( A => n1941, B => n3073, C => n870, D => n3074, Z => 
                           n4195);
   U4190 : AO4 port map( A => n1942, B => n3075, C => n871, D => n3076, Z => 
                           n4194);
   U4191 : AO4 port map( A => n1943, B => n3077, C => n872, D => n3078, Z => 
                           n4193);
   U4192 : MUX21L port map( A => n1045, B => n4197, S => CE_I, Z => n4553);
   U4193 : NR2 port map( A => n4198, B => n4199, Z => n4197);
   U4194 : ND4 port map( A => n4200, B => n4201, C => n4202, D => n4203, Z => 
                           n4199);
   U4195 : NR4 port map( A => n4204, B => n4205, C => n4206, D => n4207, Z => 
                           n4203);
   U4196 : AO4 port map( A => n1944, B => n2983, C => n873, D => n2984, Z => 
                           n4207);
   U4197 : AO4 port map( A => n1945, B => n2985, C => n874, D => n2986, Z => 
                           n4206);
   U4198 : AO4 port map( A => n1946, B => n2987, C => n875, D => n2988, Z => 
                           n4205);
   U4199 : AO4 port map( A => n1947, B => n2989, C => n876, D => n2990, Z => 
                           n4204);
   U4200 : NR4 port map( A => n4208, B => n4209, C => n4210, D => n4211, Z => 
                           n4202);
   U4201 : AO4 port map( A => n1948, B => n2995, C => n877, D => n2996, Z => 
                           n4211);
   U4202 : AO4 port map( A => n1949, B => n2997, C => n878, D => n2998, Z => 
                           n4210);
   U4203 : AO4 port map( A => n1950, B => n2999, C => n879, D => n3000, Z => 
                           n4209);
   U4204 : AO4 port map( A => n1951, B => n3001, C => n880, D => n3002, Z => 
                           n4208);
   U4205 : NR4 port map( A => n4212, B => n4213, C => n4214, D => n4215, Z => 
                           n4201);
   U4206 : AO4 port map( A => n1952, B => n3007, C => n881, D => n3008, Z => 
                           n4215);
   U4207 : AO4 port map( A => n1953, B => n3009, C => n882, D => n3010, Z => 
                           n4214);
   U4208 : AO4 port map( A => n1954, B => n3011, C => n883, D => n3012, Z => 
                           n4213);
   U4209 : AO4 port map( A => n1955, B => n3013, C => n884, D => n3014, Z => 
                           n4212);
   U4210 : NR4 port map( A => n4216, B => n4217, C => n4218, D => n4219, Z => 
                           n4200);
   U4211 : AO4 port map( A => n1956, B => n3019, C => n885, D => n3020, Z => 
                           n4219);
   U4212 : AO4 port map( A => n1957, B => n3021, C => n886, D => n3022, Z => 
                           n4218);
   U4213 : AO4 port map( A => n1958, B => n3023, C => n887, D => n3024, Z => 
                           n4217);
   U4214 : AO4 port map( A => n1959, B => n3025, C => n888, D => n3026, Z => 
                           n4216);
   U4215 : ND4 port map( A => n4220, B => n4221, C => n4222, D => n4223, Z => 
                           n4198);
   U4216 : NR4 port map( A => n4224, B => n4225, C => n4226, D => n4227, Z => 
                           n4223);
   U4217 : AO4 port map( A => n1960, B => n3035, C => n889, D => n3036, Z => 
                           n4227);
   U4218 : AO4 port map( A => n1961, B => n3037, C => n890, D => n3038, Z => 
                           n4226);
   U4219 : AO4 port map( A => n1962, B => n3039, C => n891, D => n3040, Z => 
                           n4225);
   U4220 : AO4 port map( A => n1963, B => n3041, C => n892, D => n3042, Z => 
                           n4224);
   U4221 : NR4 port map( A => n4228, B => n4229, C => n4230, D => n4231, Z => 
                           n4222);
   U4222 : AO4 port map( A => n1964, B => n3047, C => n893, D => n3048, Z => 
                           n4231);
   U4223 : AO4 port map( A => n1965, B => n3049, C => n894, D => n3050, Z => 
                           n4230);
   U4224 : AO4 port map( A => n1966, B => n3051, C => n895, D => n3052, Z => 
                           n4229);
   U4225 : AO4 port map( A => n1967, B => n3053, C => n896, D => n3054, Z => 
                           n4228);
   U4226 : NR4 port map( A => n4232, B => n4233, C => n4234, D => n4235, Z => 
                           n4221);
   U4227 : AO4 port map( A => n1968, B => n3059, C => n897, D => n3060, Z => 
                           n4235);
   U4228 : AO4 port map( A => n1969, B => n3061, C => n898, D => n3062, Z => 
                           n4234);
   U4229 : AO4 port map( A => n1970, B => n3063, C => n899, D => n3064, Z => 
                           n4233);
   U4230 : AO4 port map( A => n1971, B => n3065, C => n900, D => n3066, Z => 
                           n4232);
   U4231 : NR4 port map( A => n4236, B => n4237, C => n4238, D => n4239, Z => 
                           n4220);
   U4232 : AO4 port map( A => n1972, B => n3071, C => n901, D => n3072, Z => 
                           n4239);
   U4233 : AO4 port map( A => n1973, B => n3073, C => n902, D => n3074, Z => 
                           n4238);
   U4234 : AO4 port map( A => n1974, B => n3075, C => n903, D => n3076, Z => 
                           n4237);
   U4235 : AO4 port map( A => n1975, B => n3077, C => n904, D => n3078, Z => 
                           n4236);
   U4236 : MUX21L port map( A => n4459, B => n4240, S => CE_I, Z => n4552);
   U4237 : NR2 port map( A => n4241, B => n4242, Z => n4240);
   U4238 : ND4 port map( A => n4243, B => n4244, C => n4245, D => n4246, Z => 
                           n4242);
   U4239 : NR4 port map( A => n4247, B => n4248, C => n4249, D => n4250, Z => 
                           n4246);
   U4240 : AO4 port map( A => n1976, B => n2983, C => n905, D => n2984, Z => 
                           n4250);
   U4241 : AO4 port map( A => n1977, B => n2985, C => n906, D => n2986, Z => 
                           n4249);
   U4242 : AO4 port map( A => n1978, B => n2987, C => n907, D => n2988, Z => 
                           n4248);
   U4243 : AO4 port map( A => n1979, B => n2989, C => n908, D => n2990, Z => 
                           n4247);
   U4244 : NR4 port map( A => n4251, B => n4252, C => n4253, D => n4254, Z => 
                           n4245);
   U4245 : AO4 port map( A => n1980, B => n2995, C => n909, D => n2996, Z => 
                           n4254);
   U4246 : AO4 port map( A => n1981, B => n2997, C => n910, D => n2998, Z => 
                           n4253);
   U4247 : AO4 port map( A => n1982, B => n2999, C => n911, D => n3000, Z => 
                           n4252);
   U4248 : AO4 port map( A => n1983, B => n3001, C => n912, D => n3002, Z => 
                           n4251);
   U4249 : AO4 port map( A => n4255, B => n4256, C => n4257, D => n4258, Z => 
                           n4244);
   U4250 : AO4 port map( A => n1984, B => n3007, C => n913, D => n3008, Z => 
                           n4258);
   U4251 : AO4 port map( A => n1985, B => n3009, C => n914, D => n3010, Z => 
                           n4257);
   U4252 : AO4 port map( A => n1986, B => n3011, C => n915, D => n3012, Z => 
                           n4256);
   U4253 : AO4 port map( A => n1987, B => n3013, C => n916, D => n3014, Z => 
                           n4255);
   U4254 : NR4 port map( A => n4259, B => n4260, C => n4261, D => n4262, Z => 
                           n4243);
   U4255 : AO4 port map( A => n1988, B => n3019, C => n917, D => n3020, Z => 
                           n4262);
   U4256 : AO4 port map( A => n1989, B => n3021, C => n918, D => n3022, Z => 
                           n4261);
   U4257 : AO4 port map( A => n1990, B => n3023, C => n919, D => n3024, Z => 
                           n4260);
   U4258 : AO4 port map( A => n1991, B => n3025, C => n920, D => n3026, Z => 
                           n4259);
   U4259 : ND4 port map( A => n4263, B => n4264, C => n4265, D => n4266, Z => 
                           n4241);
   U4260 : NR4 port map( A => n4267, B => n4268, C => n4269, D => n4270, Z => 
                           n4266);
   U4261 : AO4 port map( A => n1992, B => n3035, C => n921, D => n3036, Z => 
                           n4270);
   U4262 : AO4 port map( A => n1993, B => n3037, C => n922, D => n3038, Z => 
                           n4269);
   U4263 : AO4 port map( A => n1994, B => n3039, C => n923, D => n3040, Z => 
                           n4268);
   U4264 : AO4 port map( A => n1995, B => n3041, C => n924, D => n3042, Z => 
                           n4267);
   U4265 : NR4 port map( A => n4271, B => n4272, C => n4273, D => n4274, Z => 
                           n4265);
   U4266 : AO4 port map( A => n1996, B => n3047, C => n925, D => n3048, Z => 
                           n4274);
   U4267 : AO4 port map( A => n1997, B => n3049, C => n926, D => n3050, Z => 
                           n4273);
   U4268 : AO4 port map( A => n1998, B => n3051, C => n927, D => n3052, Z => 
                           n4272);
   U4269 : AO4 port map( A => n1999, B => n3053, C => n928, D => n3054, Z => 
                           n4271);
   U4270 : NR4 port map( A => n4275, B => n4276, C => n4277, D => n4278, Z => 
                           n4264);
   U4271 : AO4 port map( A => n2000, B => n3059, C => n929, D => n3060, Z => 
                           n4278);
   U4272 : AO4 port map( A => n2001, B => n3061, C => n930, D => n3062, Z => 
                           n4277);
   U4273 : AO4 port map( A => n2002, B => n3063, C => n931, D => n3064, Z => 
                           n4276);
   U4274 : AO4 port map( A => n2003, B => n3065, C => n932, D => n3066, Z => 
                           n4275);
   U4275 : NR4 port map( A => n4279, B => n4280, C => n4281, D => n4282, Z => 
                           n4263);
   U4276 : AO4 port map( A => n2004, B => n3071, C => n933, D => n3072, Z => 
                           n4282);
   U4277 : AO4 port map( A => n2005, B => n3073, C => n934, D => n3074, Z => 
                           n4281);
   U4278 : AO4 port map( A => n2006, B => n3075, C => n935, D => n3076, Z => 
                           n4280);
   U4279 : AO4 port map( A => n2007, B => n3077, C => n936, D => n3078, Z => 
                           n4279);
   U4280 : MUX21L port map( A => n1058, B => n4283, S => CE_I, Z => n4551);
   U4281 : NR2 port map( A => n4284, B => n4285, Z => n4283);
   U4282 : ND4 port map( A => n4286, B => n4287, C => n4288, D => n4289, Z => 
                           n4285);
   U4283 : NR4 port map( A => n4290, B => n4291, C => n4292, D => n4293, Z => 
                           n4289);
   U4284 : AO4 port map( A => n2008, B => n2983, C => n937, D => n2984, Z => 
                           n4293);
   U4285 : AO4 port map( A => n2009, B => n2985, C => n938, D => n2986, Z => 
                           n4292);
   U4286 : AO4 port map( A => n2010, B => n2987, C => n939, D => n2988, Z => 
                           n4291);
   U4287 : AO4 port map( A => n2011, B => n2989, C => n940, D => n2990, Z => 
                           n4290);
   U4288 : NR4 port map( A => n4294, B => n4295, C => n4296, D => n4297, Z => 
                           n4288);
   U4289 : AO4 port map( A => n2012, B => n2995, C => n941, D => n2996, Z => 
                           n4297);
   U4290 : AO4 port map( A => n2013, B => n2997, C => n942, D => n2998, Z => 
                           n4296);
   U4291 : AO4 port map( A => n2014, B => n2999, C => n943, D => n3000, Z => 
                           n4295);
   U4292 : AO4 port map( A => n2015, B => n3001, C => n944, D => n3002, Z => 
                           n4294);
   U4293 : NR4 port map( A => n4298, B => n4299, C => n4300, D => n4301, Z => 
                           n4287);
   U4294 : AO4 port map( A => n2016, B => n3007, C => n945, D => n3008, Z => 
                           n4301);
   U4295 : AO4 port map( A => n2017, B => n3009, C => n946, D => n3010, Z => 
                           n4300);
   U4296 : AO4 port map( A => n2018, B => n3011, C => n947, D => n3012, Z => 
                           n4299);
   U4297 : AO4 port map( A => n2019, B => n3013, C => n948, D => n3014, Z => 
                           n4298);
   U4298 : NR4 port map( A => n4302, B => n4303, C => n4304, D => n4305, Z => 
                           n4286);
   U4299 : AO4 port map( A => n2020, B => n3019, C => n949, D => n3020, Z => 
                           n4305);
   U4300 : AO4 port map( A => n2021, B => n3021, C => n950, D => n3022, Z => 
                           n4304);
   U4301 : AO4 port map( A => n2022, B => n3023, C => n951, D => n3024, Z => 
                           n4303);
   U4302 : AO4 port map( A => n2023, B => n3025, C => n952, D => n3026, Z => 
                           n4302);
   U4303 : ND4 port map( A => n4306, B => n4307, C => n4308, D => n4309, Z => 
                           n4284);
   U4304 : NR4 port map( A => n4310, B => n4311, C => n4312, D => n4313, Z => 
                           n4309);
   U4305 : AO4 port map( A => n2024, B => n3035, C => n953, D => n3036, Z => 
                           n4313);
   U4306 : AO4 port map( A => n2025, B => n3037, C => n954, D => n3038, Z => 
                           n4312);
   U4307 : AO4 port map( A => n2026, B => n3039, C => n955, D => n3040, Z => 
                           n4311);
   U4308 : AO4 port map( A => n2027, B => n3041, C => n956, D => n3042, Z => 
                           n4310);
   U4309 : NR4 port map( A => n4314, B => n4315, C => n4316, D => n4317, Z => 
                           n4308);
   U4310 : AO4 port map( A => n2028, B => n3047, C => n957, D => n3048, Z => 
                           n4317);
   U4311 : AO4 port map( A => n2029, B => n3049, C => n958, D => n3050, Z => 
                           n4316);
   U4312 : AO4 port map( A => n2030, B => n3051, C => n959, D => n3052, Z => 
                           n4315);
   U4313 : AO4 port map( A => n2031, B => n3053, C => n960, D => n3054, Z => 
                           n4314);
   U4314 : NR4 port map( A => n4318, B => n4319, C => n4320, D => n4321, Z => 
                           n4307);
   U4315 : AO4 port map( A => n2032, B => n3059, C => n961, D => n3060, Z => 
                           n4321);
   U4316 : AO4 port map( A => n2033, B => n3061, C => n962, D => n3062, Z => 
                           n4320);
   U4317 : AO4 port map( A => n2034, B => n3063, C => n963, D => n3064, Z => 
                           n4319);
   U4318 : AO4 port map( A => n2035, B => n3065, C => n964, D => n3066, Z => 
                           n4318);
   U4319 : NR4 port map( A => n4322, B => n4323, C => n4324, D => n4325, Z => 
                           n4306);
   U4320 : AO4 port map( A => n2036, B => n3071, C => n965, D => n3072, Z => 
                           n4325);
   U4321 : AO4 port map( A => n2037, B => n3073, C => n966, D => n3074, Z => 
                           n4324);
   U4322 : AO4 port map( A => n2038, B => n3075, C => n967, D => n3076, Z => 
                           n4323);
   U4323 : AO4 port map( A => n2039, B => n3077, C => n968, D => n3078, Z => 
                           n4322);
   U4324 : MUX21L port map( A => n1067, B => n4326, S => CE_I, Z => n4550);
   U4325 : NR2 port map( A => n4327, B => n4328, Z => n4326);
   U4326 : ND4 port map( A => n4329, B => n4330, C => n4331, D => n4332, Z => 
                           n4328);
   U4327 : NR4 port map( A => n4333, B => n4334, C => n4335, D => n4336, Z => 
                           n4332);
   U4328 : AO4 port map( A => n2040, B => n2983, C => n969, D => n2984, Z => 
                           n4336);
   U4329 : AO4 port map( A => n2041, B => n2985, C => n970, D => n2986, Z => 
                           n4335);
   U4330 : AO4 port map( A => n2042, B => n2987, C => n971, D => n2988, Z => 
                           n4334);
   U4331 : AO4 port map( A => n2043, B => n2989, C => n972, D => n2990, Z => 
                           n4333);
   U4332 : NR4 port map( A => n4337, B => n4338, C => n4339, D => n4340, Z => 
                           n4331);
   U4333 : AO4 port map( A => n2044, B => n2995, C => n973, D => n2996, Z => 
                           n4340);
   U4334 : AO4 port map( A => n2045, B => n2997, C => n974, D => n2998, Z => 
                           n4339);
   U4335 : AO4 port map( A => n2046, B => n2999, C => n975, D => n3000, Z => 
                           n4338);
   U4336 : AO4 port map( A => n2047, B => n3001, C => n976, D => n3002, Z => 
                           n4337);
   U4337 : NR4 port map( A => n4341, B => n4342, C => n4343, D => n4344, Z => 
                           n4330);
   U4338 : AO4 port map( A => n2048, B => n3007, C => n977, D => n3008, Z => 
                           n4344);
   U4339 : AO4 port map( A => n2049, B => n3009, C => n978, D => n3010, Z => 
                           n4343);
   U4340 : AO4 port map( A => n2050, B => n3011, C => n979, D => n3012, Z => 
                           n4342);
   U4341 : AO4 port map( A => n2051, B => n3013, C => n980, D => n3014, Z => 
                           n4341);
   U4342 : NR4 port map( A => n4345, B => n4346, C => n4347, D => n4348, Z => 
                           n4329);
   U4343 : AO4 port map( A => n2052, B => n3019, C => n981, D => n3020, Z => 
                           n4348);
   U4344 : AO4 port map( A => n2053, B => n3021, C => n982, D => n3022, Z => 
                           n4347);
   U4345 : AO4 port map( A => n2054, B => n3023, C => n983, D => n3024, Z => 
                           n4346);
   U4346 : AO4 port map( A => n2055, B => n3025, C => n984, D => n3026, Z => 
                           n4345);
   U4347 : ND4 port map( A => n4349, B => n4350, C => n4351, D => n4352, Z => 
                           n4327);
   U4348 : NR4 port map( A => n4353, B => n4354, C => n4355, D => n4356, Z => 
                           n4352);
   U4349 : AO4 port map( A => n2056, B => n3035, C => n985, D => n3036, Z => 
                           n4356);
   U4350 : AO4 port map( A => n2057, B => n3037, C => n986, D => n3038, Z => 
                           n4355);
   U4351 : AO4 port map( A => n2058, B => n3039, C => n987, D => n3040, Z => 
                           n4354);
   U4352 : AO4 port map( A => n2059, B => n3041, C => n988, D => n3042, Z => 
                           n4353);
   U4353 : NR4 port map( A => n4357, B => n4358, C => n4359, D => n4360, Z => 
                           n4351);
   U4354 : AO4 port map( A => n2060, B => n3047, C => n989, D => n3048, Z => 
                           n4360);
   U4355 : AO4 port map( A => n2061, B => n3049, C => n990, D => n3050, Z => 
                           n4359);
   U4356 : AO4 port map( A => n2062, B => n3051, C => n991, D => n3052, Z => 
                           n4358);
   U4357 : AO4 port map( A => n2063, B => n3053, C => n992, D => n3054, Z => 
                           n4357);
   U4358 : NR4 port map( A => n4361, B => n4362, C => n4363, D => n4364, Z => 
                           n4350);
   U4359 : AO4 port map( A => n2064, B => n3059, C => n993, D => n3060, Z => 
                           n4364);
   U4360 : AO4 port map( A => n2065, B => n3061, C => n994, D => n3062, Z => 
                           n4363);
   U4361 : AO4 port map( A => n2066, B => n3063, C => n995, D => n3064, Z => 
                           n4362);
   U4362 : AO4 port map( A => n2067, B => n3065, C => n996, D => n3066, Z => 
                           n4361);
   U4363 : NR4 port map( A => n4365, B => n4366, C => n4367, D => n4368, Z => 
                           n4349);
   U4364 : AO4 port map( A => n2068, B => n3071, C => n997, D => n3072, Z => 
                           n4368);
   U4365 : AO4 port map( A => n2069, B => n3073, C => n998, D => n3074, Z => 
                           n4367);
   U4366 : AO4 port map( A => n2070, B => n3075, C => n999, D => n3076, Z => 
                           n4366);
   U4367 : AO4 port map( A => n2071, B => n3077, C => n1000, D => n3078, Z => 
                           n4365);
   U4368 : MUX21L port map( A => n1046, B => n4369, S => CE_I, Z => n4549);
   U4369 : NR2 port map( A => n4370, B => n4371, Z => n4369);
   U4370 : ND4 port map( A => n4372, B => n4373, C => n4374, D => n4375, Z => 
                           n4371);
   U4371 : NR4 port map( A => n4376, B => n4377, C => n4378, D => n4379, Z => 
                           n4375);
   U4372 : AO4 port map( A => n2072, B => n2983, C => n1001, D => n2984, Z => 
                           n4379);
   U4373 : ND2 port map( A => n4380, B => n4381, Z => n2984);
   U4374 : ND2 port map( A => n4380, B => n4382, Z => n2983);
   U4375 : AO4 port map( A => n2073, B => n2985, C => n1002, D => n2986, Z => 
                           n4378);
   U4376 : ND2 port map( A => n4380, B => n4383, Z => n2986);
   U4377 : ND2 port map( A => n4380, B => n4384, Z => n2985);
   U4378 : AN2 port map( A => n4385, B => n4386, Z => n4380);
   U4379 : AO4 port map( A => n2074, B => n2987, C => n1003, D => n2988, Z => 
                           n4377);
   U4380 : ND2 port map( A => n4387, B => n4381, Z => n2988);
   U4381 : ND2 port map( A => n4387, B => n4382, Z => n2987);
   U4382 : AO4 port map( A => n2075, B => n2989, C => n1004, D => n2990, Z => 
                           n4376);
   U4383 : ND2 port map( A => n4387, B => n4383, Z => n2990);
   U4384 : ND2 port map( A => n4387, B => n4384, Z => n2989);
   U4385 : AN2 port map( A => n4385, B => n4388, Z => n4387);
   U4386 : NR4 port map( A => n4389, B => n4390, C => n4391, D => n4392, Z => 
                           n4374);
   U4387 : AO4 port map( A => n2076, B => n2995, C => n1005, D => n2996, Z => 
                           n4392);
   U4388 : ND2 port map( A => n4393, B => n4381, Z => n2996);
   U4389 : ND2 port map( A => n4393, B => n4382, Z => n2995);
   U4390 : AO4 port map( A => n2077, B => n2997, C => n1006, D => n2998, Z => 
                           n4391);
   U4391 : ND2 port map( A => n4393, B => n4383, Z => n2998);
   U4392 : ND2 port map( A => n4393, B => n4384, Z => n2997);
   U4393 : AN2 port map( A => n4385, B => n4394, Z => n4393);
   U4394 : AO4 port map( A => n2078, B => n2999, C => n1007, D => n3000, Z => 
                           n4390);
   U4395 : ND2 port map( A => n4395, B => n4381, Z => n3000);
   U4396 : ND2 port map( A => n4395, B => n4382, Z => n2999);
   U4397 : AO4 port map( A => n2079, B => n3001, C => n1008, D => n3002, Z => 
                           n4389);
   U4398 : ND2 port map( A => n4395, B => n4383, Z => n3002);
   U4399 : ND2 port map( A => n4395, B => n4384, Z => n3001);
   U4400 : AN2 port map( A => n4385, B => n4396, Z => n4395);
   U4401 : NR2 port map( A => n4397, B => n4398, Z => n4385);
   U4402 : NR4 port map( A => n4399, B => n4400, C => n4401, D => n4402, Z => 
                           n4373);
   U4403 : AO4 port map( A => n2080, B => n3007, C => n1009, D => n3008, Z => 
                           n4402);
   U4404 : ND2 port map( A => n4403, B => n4381, Z => n3008);
   U4405 : ND2 port map( A => n4403, B => n4382, Z => n3007);
   U4406 : AO4 port map( A => n2081, B => n3009, C => n1010, D => n3010, Z => 
                           n4401);
   U4407 : ND2 port map( A => n4403, B => n4383, Z => n3010);
   U4408 : ND2 port map( A => n4403, B => n4384, Z => n3009);
   U4409 : AN2 port map( A => n4404, B => n4386, Z => n4403);
   U4410 : AO4 port map( A => n2082, B => n3011, C => n1011, D => n3012, Z => 
                           n4400);
   U4411 : ND2 port map( A => n4405, B => n4381, Z => n3012);
   U4412 : ND2 port map( A => n4405, B => n4382, Z => n3011);
   U4413 : AO4 port map( A => n2083, B => n3013, C => n1012, D => n3014, Z => 
                           n4399);
   U4414 : ND2 port map( A => n4405, B => n4383, Z => n3014);
   U4415 : ND2 port map( A => n4405, B => n4384, Z => n3013);
   U4416 : AN2 port map( A => n4404, B => n4388, Z => n4405);
   U4417 : NR4 port map( A => n4406, B => n4407, C => n4408, D => n4409, Z => 
                           n4372);
   U4418 : AO4 port map( A => n2084, B => n3019, C => n1013, D => n3020, Z => 
                           n4409);
   U4419 : ND2 port map( A => n4410, B => n4381, Z => n3020);
   U4420 : ND2 port map( A => n4410, B => n4382, Z => n3019);
   U4421 : AO4 port map( A => n2085, B => n3021, C => n1014, D => n3022, Z => 
                           n4408);
   U4422 : ND2 port map( A => n4410, B => n4383, Z => n3022);
   U4423 : ND2 port map( A => n4410, B => n4384, Z => n3021);
   U4424 : AN2 port map( A => n4404, B => n4394, Z => n4410);
   U4425 : AO4 port map( A => n2086, B => n3023, C => n1015, D => n3024, Z => 
                           n4407);
   U4426 : ND2 port map( A => n4411, B => n4381, Z => n3024);
   U4427 : ND2 port map( A => n4411, B => n4382, Z => n3023);
   U4428 : AO4 port map( A => n2087, B => n3025, C => n1016, D => n3026, Z => 
                           n4406);
   U4429 : ND2 port map( A => n4411, B => n4383, Z => n3026);
   U4430 : ND2 port map( A => n4411, B => n4384, Z => n3025);
   U4431 : AN2 port map( A => n4404, B => n4396, Z => n4411);
   U4432 : NR2 port map( A => n4398, B => n4412, Z => n4404);
   U4433 : ND4 port map( A => n4413, B => n4414, C => n4415, D => n4416, Z => 
                           n4370);
   U4434 : NR4 port map( A => n4417, B => n4418, C => n4419, D => n4420, Z => 
                           n4416);
   U4435 : AO4 port map( A => n2088, B => n3035, C => n1017, D => n3036, Z => 
                           n4420);
   U4436 : ND2 port map( A => n4421, B => n4381, Z => n3036);
   U4437 : ND2 port map( A => n4421, B => n4382, Z => n3035);
   U4438 : AO4 port map( A => n2089, B => n3037, C => n1018, D => n3038, Z => 
                           n4419);
   U4439 : ND2 port map( A => n4421, B => n4383, Z => n3038);
   U4440 : ND2 port map( A => n4421, B => n4384, Z => n3037);
   U4441 : AN2 port map( A => n4386, B => n4422, Z => n4421);
   U4442 : AO4 port map( A => n2090, B => n3039, C => n1019, D => n3040, Z => 
                           n4418);
   U4443 : ND2 port map( A => n4381, B => n4423, Z => n3040);
   U4444 : ND2 port map( A => n4382, B => n4423, Z => n3039);
   U4445 : AO4 port map( A => n2091, B => n3041, C => n1020, D => n3042, Z => 
                           n4417);
   U4446 : ND2 port map( A => n4423, B => n4383, Z => n3042);
   U4447 : ND2 port map( A => n4384, B => n4423, Z => n3041);
   U4448 : AN2 port map( A => n4422, B => n4388, Z => n4423);
   U4449 : NR4 port map( A => n4424, B => n4425, C => n4426, D => n4427, Z => 
                           n4415);
   U4450 : AO4 port map( A => n2092, B => n3047, C => n1021, D => n3048, Z => 
                           n4427);
   U4451 : ND2 port map( A => n4428, B => n4381, Z => n3048);
   U4452 : ND2 port map( A => n4428, B => n4382, Z => n3047);
   U4453 : AO4 port map( A => n2093, B => n3049, C => n1022, D => n3050, Z => 
                           n4426);
   U4454 : ND2 port map( A => n4428, B => n4383, Z => n3050);
   U4455 : ND2 port map( A => n4428, B => n4384, Z => n3049);
   U4456 : AN2 port map( A => n4394, B => n4422, Z => n4428);
   U4457 : AO4 port map( A => n2094, B => n3051, C => n1023, D => n3052, Z => 
                           n4425);
   U4458 : ND2 port map( A => n4429, B => n4381, Z => n3052);
   U4459 : ND2 port map( A => n4429, B => n4382, Z => n3051);
   U4460 : AO4 port map( A => n2095, B => n3053, C => n1024, D => n3054, Z => 
                           n4424);
   U4461 : ND2 port map( A => n4429, B => n4383, Z => n3054);
   U4462 : ND2 port map( A => n4429, B => n4384, Z => n3053);
   U4463 : AN2 port map( A => n4396, B => n4422, Z => n4429);
   U4464 : NR2 port map( A => n4397, B => n4430, Z => n4422);
   U4465 : NR4 port map( A => n4431, B => n4432, C => n4433, D => n4434, Z => 
                           n4414);
   U4466 : AO4 port map( A => n2096, B => n3059, C => n1025, D => n3060, Z => 
                           n4434);
   U4467 : ND2 port map( A => n4435, B => n4381, Z => n3060);
   U4468 : ND2 port map( A => n4435, B => n4382, Z => n3059);
   U4469 : AO4 port map( A => n2097, B => n3061, C => n1026, D => n3062, Z => 
                           n4433);
   U4470 : ND2 port map( A => n4435, B => n4383, Z => n3062);
   U4471 : ND2 port map( A => n4435, B => n4384, Z => n3061);
   U4472 : AN2 port map( A => n4436, B => n4386, Z => n4435);
   U4473 : NR2 port map( A => n4437, B => n4438, Z => n4386);
   U4474 : AO4 port map( A => n2098, B => n3063, C => n1027, D => n3064, Z => 
                           n4432);
   U4475 : ND2 port map( A => n4439, B => n4381, Z => n3064);
   U4476 : ND2 port map( A => n4439, B => n4382, Z => n3063);
   U4477 : AO4 port map( A => n2099, B => n3065, C => n1028, D => n3066, Z => 
                           n4431);
   U4478 : ND2 port map( A => n4439, B => n4383, Z => n3066);
   U4479 : ND2 port map( A => n4439, B => n4384, Z => n3065);
   U4480 : AN2 port map( A => n4436, B => n4388, Z => n4439);
   U4481 : NR2 port map( A => n4437, B => n4440, Z => n4388);
   U4482 : NR4 port map( A => n4441, B => n4442, C => n4443, D => n4444, Z => 
                           n4413);
   U4483 : AO4 port map( A => n2100, B => n3071, C => n1029, D => n3072, Z => 
                           n4444);
   U4484 : ND2 port map( A => n4445, B => n4381, Z => n3072);
   U4485 : ND2 port map( A => n4445, B => n4382, Z => n3071);
   U4486 : AO4 port map( A => n2101, B => n3073, C => n1030, D => n3074, Z => 
                           n4443);
   U4487 : ND2 port map( A => n4445, B => n4383, Z => n3074);
   U4488 : ND2 port map( A => n4445, B => n4384, Z => n3073);
   U4489 : AN2 port map( A => n4436, B => n4394, Z => n4445);
   U4490 : NR2 port map( A => n4438, B => n4446, Z => n4394);
   U4491 : AO4 port map( A => n2102, B => n3075, C => n1031, D => n3076, Z => 
                           n4442);
   U4492 : ND2 port map( A => n4447, B => n4381, Z => n3076);
   U4493 : NR2 port map( A => n4448, B => n4449, Z => n4381);
   U4494 : ND2 port map( A => n4447, B => n4382, Z => n3075);
   U4495 : NR2 port map( A => n4450, B => n4449, Z => n4382);
   U4496 : IV port map( A => n4451, Z => n4449);
   U4497 : AO4 port map( A => n2103, B => n3077, C => n1032, D => n3078, Z => 
                           n4441);
   U4498 : ND2 port map( A => n4447, B => n4383, Z => n3078);
   U4499 : NR2 port map( A => n4451, B => n4448, Z => n4383);
   U4500 : IV port map( A => n4450, Z => n4448);
   U4501 : ND2 port map( A => n4447, B => n4384, Z => n3077);
   U4502 : NR2 port map( A => n4450, B => n4451, Z => n4384);
   U4503 : MUX21L port map( A => n1033, B => KEY_NUMB_I(1), S => GET_KEY_I, Z 
                           => n4451);
   U4504 : MUX21L port map( A => n1, B => KEY_NUMB_I(0), S => GET_KEY_I, Z => 
                           n4450);
   U4505 : AN2 port map( A => n4436, B => n4396, Z => n4447);
   U4506 : NR2 port map( A => n4440, B => n4446, Z => n4396);
   U4507 : IV port map( A => n4437, Z => n4446);
   U4508 : MUX21L port map( A => n1044, B => KEY_NUMB_I(3), S => GET_KEY_I, Z 
                           => n4437);
   U4509 : IV port map( A => n4438, Z => n4440);
   U4510 : MUX21L port map( A => n6647, B => n4452, S => GET_KEY_I, Z => n4438)
                           ;
   U4511 : IV port map( A => KEY_NUMB_I(2), Z => n4452);
   U4512 : NR2 port map( A => n4430, B => n4412, Z => n4436);
   U4513 : IV port map( A => n4397, Z => n4412);
   U4514 : MUX21L port map( A => n1037, B => KEY_NUMB_I(4), S => GET_KEY_I, Z 
                           => n4397);
   U4515 : IV port map( A => n4398, Z => n4430);
   U4516 : MUX21L port map( A => n6644, B => n4453, S => GET_KEY_I, Z => n4398)
                           ;
   U4517 : IV port map( A => KEY_NUMB_I(5), Z => n4453);
   U4518 : NR2 port map( A => n1045, B => n1034, Z => KEY_EXP_O(9));
   U4519 : NR2 port map( A => n1046, B => n1034, Z => KEY_EXP_O(8));
   U4520 : NR2 port map( A => n4454, B => n1034, Z => KEY_EXP_O(7));
   U4521 : NR2 port map( A => n4457, B => n1034, Z => KEY_EXP_O(6));
   U4522 : NR2 port map( A => n1047, B => n1034, Z => KEY_EXP_O(5));
   U4523 : NR2 port map( A => n1048, B => n1034, Z => KEY_EXP_O(4));
   U4524 : NR2 port map( A => n1049, B => n1034, Z => KEY_EXP_O(3));
   U4525 : NR2 port map( A => n1050, B => n1034, Z => KEY_EXP_O(31));
   U4526 : NR2 port map( A => n1051, B => n1034, Z => KEY_EXP_O(30));
   U4527 : NR2 port map( A => n1052, B => n1034, Z => KEY_EXP_O(2));
   U4528 : NR2 port map( A => n1053, B => n1034, Z => KEY_EXP_O(29));
   U4529 : NR2 port map( A => n1054, B => n1034, Z => KEY_EXP_O(28));
   U4530 : NR2 port map( A => n1055, B => n1034, Z => KEY_EXP_O(27));
   U4531 : NR2 port map( A => n1056, B => n1034, Z => KEY_EXP_O(26));
   U4532 : NR2 port map( A => n1057, B => n1034, Z => KEY_EXP_O(25));
   U4533 : NR2 port map( A => n1058, B => n1034, Z => KEY_EXP_O(24));
   U4534 : NR2 port map( A => n1059, B => n1034, Z => KEY_EXP_O(23));
   U4535 : NR2 port map( A => n1060, B => n1034, Z => KEY_EXP_O(22));
   U4536 : NR2 port map( A => n1061, B => n1034, Z => KEY_EXP_O(21));
   U4537 : NR2 port map( A => n1062, B => n1034, Z => KEY_EXP_O(20));
   U4538 : NR2 port map( A => n1063, B => n1034, Z => KEY_EXP_O(1));
   U4539 : NR2 port map( A => n1064, B => n1034, Z => KEY_EXP_O(19));
   U4540 : NR2 port map( A => n1065, B => n1034, Z => KEY_EXP_O(18));
   U4541 : NR2 port map( A => n1066, B => n1034, Z => KEY_EXP_O(17));
   U4542 : NR2 port map( A => n1067, B => n1034, Z => KEY_EXP_O(16));
   U4543 : NR2 port map( A => n1068, B => n1034, Z => KEY_EXP_O(15));
   U4544 : NR2 port map( A => n1069, B => n1034, Z => KEY_EXP_O(14));
   U4545 : NR2 port map( A => n1070, B => n1034, Z => KEY_EXP_O(13));
   U4546 : NR2 port map( A => n1071, B => n1034, Z => KEY_EXP_O(12));
   U4547 : NR2 port map( A => n1072, B => n1034, Z => KEY_EXP_O(11));
   U4548 : NR2 port map( A => n1073, B => n1034, Z => KEY_EXP_O(10));
   U4549 : NR2 port map( A => n4459, B => n1034, Z => KEY_EXP_O(0));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_aes_dec_KEY_SIZE2.all;

entity aes_dec_KEY_SIZE2 is

   port( DATA_I : in std_logic_vector (7 downto 0);  VALID_DATA_I : in 
         std_logic;  KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, 
         RESET_I, CLK_I, CE_I : in std_logic;  KEY_READY_O, VALID_O : out 
         std_logic;  DATA_O : out std_logic_vector (7 downto 0));

end aes_dec_KEY_SIZE2;

architecture SYN_Behavioral of aes_dec_KEY_SIZE2 is

   component NR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component IV
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO7
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AN2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component ND3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21L
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AO3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21H
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component EN
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EO
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX31L
      port( D0, D1, D2, A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EON1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AN4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component key_expansion
      port( KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, CLK_I, 
            RESET_I, CE_I : in std_logic;  DONE_O : out std_logic;  GET_KEY_I :
            in std_logic;  KEY_NUMB_I : in std_logic_vector (5 downto 0);  
            KEY_EXP_O : out std_logic_vector (31 downto 0));
   end component;
   
   component FD1
      port( D, CP : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_O_7_port, DATA_O_6_port, DATA_O_5_port, DATA_O_4_port, 
      DATA_O_3_port, DATA_O_2_port, DATA_O_1_port, DATA_O_0_port, GET_KEY, 
      v_INV_KEY_NUMB_5_port, v_INV_KEY_NUMB_4_port, v_INV_KEY_NUMB_3_port, 
      v_INV_KEY_NUMB_2_port, v_KEY_COLUMN_31_port, v_KEY_COLUMN_30_port, 
      v_KEY_COLUMN_29_port, v_KEY_COLUMN_28_port, v_KEY_COLUMN_27_port, 
      v_KEY_COLUMN_26_port, v_KEY_COLUMN_25_port, v_KEY_COLUMN_24_port, 
      v_KEY_COLUMN_23_port, v_KEY_COLUMN_22_port, v_KEY_COLUMN_21_port, 
      v_KEY_COLUMN_20_port, v_KEY_COLUMN_19_port, v_KEY_COLUMN_18_port, 
      v_KEY_COLUMN_17_port, v_KEY_COLUMN_16_port, v_KEY_COLUMN_15_port, 
      v_KEY_COLUMN_14_port, v_KEY_COLUMN_13_port, v_KEY_COLUMN_12_port, 
      v_KEY_COLUMN_11_port, v_KEY_COLUMN_10_port, v_KEY_COLUMN_9_port, 
      v_KEY_COLUMN_8_port, v_KEY_COLUMN_7_port, v_KEY_COLUMN_6_port, 
      v_KEY_COLUMN_5_port, v_KEY_COLUMN_4_port, v_KEY_COLUMN_3_port, 
      v_KEY_COLUMN_2_port, v_KEY_COLUMN_1_port, v_KEY_COLUMN_0_port, 
      v_KEY_NUMB_1_port, v_KEY_NUMB_0_port, v_CNT4_1_port, v_CNT4_0_port, 
      v_DATA_COLUMN_31_port, v_DATA_COLUMN_30_port, v_DATA_COLUMN_29_port, 
      v_DATA_COLUMN_28_port, v_DATA_COLUMN_27_port, v_DATA_COLUMN_26_port, 
      v_DATA_COLUMN_25_port, v_DATA_COLUMN_24_port, v_DATA_COLUMN_23_port, 
      v_DATA_COLUMN_22_port, v_DATA_COLUMN_21_port, v_DATA_COLUMN_20_port, 
      v_DATA_COLUMN_19_port, v_DATA_COLUMN_18_port, v_DATA_COLUMN_17_port, 
      v_DATA_COLUMN_16_port, v_DATA_COLUMN_15_port, v_DATA_COLUMN_14_port, 
      v_DATA_COLUMN_13_port, v_DATA_COLUMN_12_port, v_DATA_COLUMN_11_port, 
      v_DATA_COLUMN_10_port, v_DATA_COLUMN_9_port, v_DATA_COLUMN_8_port, 
      v_DATA_COLUMN_7_port, v_DATA_COLUMN_6_port, v_DATA_COLUMN_5_port, 
      v_DATA_COLUMN_4_port, v_DATA_COLUMN_3_port, v_DATA_COLUMN_2_port, 
      v_DATA_COLUMN_1_port, v_DATA_COLUMN_0_port, v_CALCULATION_CNTR_7_port, 
      v_CALCULATION_CNTR_6_port, v_CALCULATION_CNTR_5_port, 
      v_CALCULATION_CNTR_4_port, v_CALCULATION_CNTR_3_port, 
      v_CALCULATION_CNTR_2_port, v_CALCULATION_CNTR_1_port, 
      v_CALCULATION_CNTR_0_port, N192, v_RAM_IN0_31_port, v_RAM_IN0_30_port, 
      v_RAM_IN0_29_port, v_RAM_IN0_28_port, v_RAM_IN0_27_port, 
      v_RAM_IN0_26_port, v_RAM_IN0_25_port, v_RAM_IN0_24_port, 
      v_RAM_IN0_23_port, v_RAM_IN0_22_port, v_RAM_IN0_21_port, 
      v_RAM_IN0_20_port, v_RAM_IN0_19_port, v_RAM_IN0_18_port, 
      v_RAM_IN0_17_port, v_RAM_IN0_16_port, v_RAM_IN0_15_port, 
      v_RAM_IN0_14_port, v_RAM_IN0_13_port, v_RAM_IN0_12_port, 
      v_RAM_IN0_11_port, v_RAM_IN0_10_port, v_RAM_IN0_9_port, v_RAM_IN0_8_port,
      v_RAM_IN0_7_port, v_RAM_IN0_6_port, v_RAM_IN0_5_port, v_RAM_IN0_4_port, 
      v_RAM_IN0_3_port, v_RAM_IN0_2_port, v_RAM_IN0_1_port, v_RAM_IN0_0_port, 
      t_STATE_RAM0_0_31_port, t_STATE_RAM0_0_29_port, t_STATE_RAM0_0_28_port, 
      t_STATE_RAM0_0_27_port, t_STATE_RAM0_0_26_port, t_STATE_RAM0_0_25_port, 
      t_STATE_RAM0_0_21_port, t_STATE_RAM0_0_20_port, t_STATE_RAM0_0_19_port, 
      t_STATE_RAM0_0_18_port, t_STATE_RAM0_0_17_port, t_STATE_RAM0_0_15_port, 
      t_STATE_RAM0_0_13_port, t_STATE_RAM0_0_12_port, t_STATE_RAM0_0_11_port, 
      t_STATE_RAM0_0_10_port, t_STATE_RAM0_0_9_port, t_STATE_RAM0_0_8_port, 
      t_STATE_RAM0_0_7_port, t_STATE_RAM0_0_5_port, t_STATE_RAM0_0_4_port, 
      t_STATE_RAM0_0_3_port, t_STATE_RAM0_0_2_port, t_STATE_RAM0_0_1_port, 
      t_STATE_RAM0_0_0_port, t_STATE_RAM0_1_31_port, t_STATE_RAM0_1_30_port, 
      t_STATE_RAM0_1_29_port, t_STATE_RAM0_1_28_port, t_STATE_RAM0_1_27_port, 
      t_STATE_RAM0_1_26_port, t_STATE_RAM0_1_25_port, t_STATE_RAM0_1_24_port, 
      t_STATE_RAM0_1_23_port, t_STATE_RAM0_1_22_port, t_STATE_RAM0_1_21_port, 
      t_STATE_RAM0_1_20_port, t_STATE_RAM0_1_19_port, t_STATE_RAM0_1_18_port, 
      t_STATE_RAM0_1_17_port, t_STATE_RAM0_1_16_port, t_STATE_RAM0_1_15_port, 
      t_STATE_RAM0_1_14_port, t_STATE_RAM0_1_13_port, t_STATE_RAM0_1_12_port, 
      t_STATE_RAM0_1_11_port, t_STATE_RAM0_1_10_port, t_STATE_RAM0_1_9_port, 
      t_STATE_RAM0_1_8_port, t_STATE_RAM0_1_7_port, t_STATE_RAM0_1_6_port, 
      t_STATE_RAM0_1_5_port, t_STATE_RAM0_1_4_port, t_STATE_RAM0_1_3_port, 
      t_STATE_RAM0_1_2_port, t_STATE_RAM0_1_1_port, t_STATE_RAM0_1_0_port, 
      t_STATE_RAM0_2_31_port, t_STATE_RAM0_2_30_port, t_STATE_RAM0_2_29_port, 
      t_STATE_RAM0_2_28_port, t_STATE_RAM0_2_27_port, t_STATE_RAM0_2_26_port, 
      t_STATE_RAM0_2_25_port, t_STATE_RAM0_2_24_port, t_STATE_RAM0_2_23_port, 
      t_STATE_RAM0_2_22_port, t_STATE_RAM0_2_21_port, t_STATE_RAM0_2_20_port, 
      t_STATE_RAM0_2_19_port, t_STATE_RAM0_2_18_port, t_STATE_RAM0_2_17_port, 
      t_STATE_RAM0_2_16_port, t_STATE_RAM0_2_15_port, t_STATE_RAM0_2_14_port, 
      t_STATE_RAM0_2_13_port, t_STATE_RAM0_2_12_port, t_STATE_RAM0_2_11_port, 
      t_STATE_RAM0_2_10_port, t_STATE_RAM0_2_9_port, t_STATE_RAM0_2_8_port, 
      t_STATE_RAM0_2_7_port, t_STATE_RAM0_2_6_port, t_STATE_RAM0_2_5_port, 
      t_STATE_RAM0_2_4_port, t_STATE_RAM0_2_3_port, t_STATE_RAM0_2_2_port, 
      t_STATE_RAM0_2_1_port, t_STATE_RAM0_2_0_port, t_STATE_RAM0_3_31_port, 
      t_STATE_RAM0_3_30_port, t_STATE_RAM0_3_29_port, t_STATE_RAM0_3_28_port, 
      t_STATE_RAM0_3_27_port, t_STATE_RAM0_3_26_port, t_STATE_RAM0_3_25_port, 
      t_STATE_RAM0_3_24_port, t_STATE_RAM0_3_23_port, t_STATE_RAM0_3_22_port, 
      t_STATE_RAM0_3_21_port, t_STATE_RAM0_3_20_port, t_STATE_RAM0_3_19_port, 
      t_STATE_RAM0_3_18_port, t_STATE_RAM0_3_17_port, t_STATE_RAM0_3_16_port, 
      t_STATE_RAM0_3_15_port, t_STATE_RAM0_3_14_port, t_STATE_RAM0_3_13_port, 
      t_STATE_RAM0_3_12_port, t_STATE_RAM0_3_11_port, t_STATE_RAM0_3_10_port, 
      t_STATE_RAM0_3_9_port, t_STATE_RAM0_3_8_port, t_STATE_RAM0_3_7_port, 
      t_STATE_RAM0_3_6_port, t_STATE_RAM0_3_5_port, t_STATE_RAM0_3_4_port, 
      t_STATE_RAM0_3_3_port, t_STATE_RAM0_3_2_port, t_STATE_RAM0_3_1_port, 
      t_STATE_RAM0_3_0_port, v_RAM_OUT0_31_port, v_RAM_OUT0_30_port, 
      v_RAM_OUT0_29_port, v_RAM_OUT0_28_port, v_RAM_OUT0_27_port, 
      v_RAM_OUT0_26_port, v_RAM_OUT0_25_port, v_RAM_OUT0_24_port, 
      v_RAM_OUT0_23_port, v_RAM_OUT0_22_port, v_RAM_OUT0_21_port, 
      v_RAM_OUT0_20_port, v_RAM_OUT0_19_port, v_RAM_OUT0_18_port, 
      v_RAM_OUT0_17_port, v_RAM_OUT0_16_port, v_RAM_OUT0_15_port, 
      v_RAM_OUT0_14_port, v_RAM_OUT0_13_port, v_RAM_OUT0_12_port, 
      v_RAM_OUT0_11_port, v_RAM_OUT0_10_port, v_RAM_OUT0_9_port, 
      v_RAM_OUT0_8_port, v_RAM_OUT0_7_port, v_RAM_OUT0_6_port, 
      v_RAM_OUT0_5_port, v_RAM_OUT0_4_port, v_RAM_OUT0_3_port, 
      v_RAM_OUT0_2_port, v_RAM_OUT0_1_port, v_RAM_OUT0_0_port, n3813, n3947, 
      n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, 
      n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, 
      n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, 
      n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, 
      n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, 
      n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, 
      n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, 
      n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, 
      n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, 
      n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, 
      n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, 
      n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, 
      n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, 
      n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, 
      n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, 
      n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, 
      n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, 
      n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, 
      n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, 
      n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, 
      n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, 
      n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, 
      n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, 
      n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, 
      n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, 
      n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, 
      n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, 
      n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, 
      n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, 
      n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, 
      n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, 
      n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, 
      n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, 
      n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, 
      n4300, n4301, n4303, n4304, n4305, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4323, n4331, n4339, n4340, n4348, n4349, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, 
      n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
      n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
      n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, 
      n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, 
      n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
      n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, 
      n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, 
      n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, 
      n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, 
      n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, 
      n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
      n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
      n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
      n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, 
      n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, 
      n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, 
      n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, 
      n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, 
      n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, 
      n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, 
      n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, 
      n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, 
      n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, 
      n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, 
      n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, 
      n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, 
      n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, 
      n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
      n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
      n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, 
      n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, 
      n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, 
      n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, 
      n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, 
      n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, 
      n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, 
      n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, 
      n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, 
      n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, 
      n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, 
      n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, 
      n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
      n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, 
      n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, 
      n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, 
      n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, 
      n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, 
      n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, 
      n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, 
      n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, 
      n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, 
      n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, 
      n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, 
      n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
      n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, 
      n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, 
      n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, 
      n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, 
      n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, 
      n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, 
      n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, 
      n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, 
      n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, 
      n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, 
      n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, 
      n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, 
      n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, 
      n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, 
      n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, 
      n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, 
      n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, 
      n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, 
      n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, 
      n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, 
      n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, 
      n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, 
      n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, 
      n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, 
      n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, 
      n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, 
      n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, 
      n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, 
      n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, 
      n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, 
      n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
      n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, 
      n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, 
      n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, 
      n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
      n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
      n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, 
      n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, 
      n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, 
      n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
      n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, 
      n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, 
      n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, 
      n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, 
      n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, 
      n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, 
      n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, 
      n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, 
      n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, 
      n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
      n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, 
      n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, 
      n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, 
      n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, 
      n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, 
      n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, 
      n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, 
      n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, 
      n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, 
      n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, 
      n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, 
      n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
      n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, 
      n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, 
      n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, 
      n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
      n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, 
      n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, 
      n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, 
      n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, 
      n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, 
      n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, 
      n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
      n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, 
      n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
      n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, 
      n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, 
      n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, 
      n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, 
      n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, 
      n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, 
      n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
      n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, 
      n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
      n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
      n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
      n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, 
      n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, 
      n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
      n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, 
      n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, 
      n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, 
      n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
      n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, 
      n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, 
      n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
      n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, 
      n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
      n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, 
      n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
      n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, 
      n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n_3112, n_3113, n_3114, n_3115, n_3116, 
      n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, 
      n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, 
      n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, 
      n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, 
      n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, 
      n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, 
      n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, 
      n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, 
      n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, 
      n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, 
      n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, 
      n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, 
      n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, 
      n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, 
      n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, 
      n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, 
      n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, 
      n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, 
      n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, 
      n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, 
      n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, 
      n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, 
      n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, 
      n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, 
      n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, 
      n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, 
      n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, 
      n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368 : 
      std_logic;

begin
   DATA_O <= ( DATA_O_7_port, DATA_O_6_port, DATA_O_5_port, DATA_O_4_port, 
      DATA_O_3_port, DATA_O_2_port, DATA_O_1_port, DATA_O_0_port );
   
   GET_KEY_reg : FD1 port map( D => N192, CP => CLK_I, Q => GET_KEY, QN => 
                           n_3112);
   v_CNT4_reg_0_inst : FD1 port map( D => n4349, CP => CLK_I, Q => 
                           v_CNT4_0_port, QN => n4418);
   v_DATA_COLUMN_reg_24_inst : FD1 port map( D => n4348, CP => CLK_I, Q => 
                           v_DATA_COLUMN_24_port, QN => n_3113);
   v_DATA_COLUMN_reg_25_inst : FD1 port map( D => n7971, CP => CLK_I, Q => 
                           v_DATA_COLUMN_25_port, QN => n_3114);
   v_DATA_COLUMN_reg_26_inst : FD1 port map( D => n7967, CP => CLK_I, Q => 
                           v_DATA_COLUMN_26_port, QN => n_3115);
   v_DATA_COLUMN_reg_27_inst : FD1 port map( D => n7963, CP => CLK_I, Q => 
                           v_DATA_COLUMN_27_port, QN => n_3116);
   v_DATA_COLUMN_reg_28_inst : FD1 port map( D => n7959, CP => CLK_I, Q => 
                           v_DATA_COLUMN_28_port, QN => n_3117);
   v_DATA_COLUMN_reg_29_inst : FD1 port map( D => n7955, CP => CLK_I, Q => 
                           v_DATA_COLUMN_29_port, QN => n_3118);
   v_DATA_COLUMN_reg_30_inst : FD1 port map( D => n7951, CP => CLK_I, Q => 
                           v_DATA_COLUMN_30_port, QN => n_3119);
   v_DATA_COLUMN_reg_31_inst : FD1 port map( D => n7947, CP => CLK_I, Q => 
                           v_DATA_COLUMN_31_port, QN => n_3120);
   v_CNT4_reg_1_inst : FD1 port map( D => n4340, CP => CLK_I, Q => 
                           v_CNT4_1_port, QN => n4370);
   v_DATA_COLUMN_reg_8_inst : FD1 port map( D => n4339, CP => CLK_I, Q => 
                           v_DATA_COLUMN_8_port, QN => n_3121);
   v_DATA_COLUMN_reg_9_inst : FD1 port map( D => n7970, CP => CLK_I, Q => 
                           v_DATA_COLUMN_9_port, QN => n_3122);
   v_DATA_COLUMN_reg_10_inst : FD1 port map( D => n7969, CP => CLK_I, Q => 
                           v_DATA_COLUMN_10_port, QN => n_3123);
   v_DATA_COLUMN_reg_11_inst : FD1 port map( D => n7965, CP => CLK_I, Q => 
                           v_DATA_COLUMN_11_port, QN => n_3124);
   v_DATA_COLUMN_reg_12_inst : FD1 port map( D => n7961, CP => CLK_I, Q => 
                           v_DATA_COLUMN_12_port, QN => n_3125);
   v_DATA_COLUMN_reg_13_inst : FD1 port map( D => n7957, CP => CLK_I, Q => 
                           v_DATA_COLUMN_13_port, QN => n_3126);
   v_DATA_COLUMN_reg_14_inst : FD1 port map( D => n7953, CP => CLK_I, Q => 
                           v_DATA_COLUMN_14_port, QN => n_3127);
   v_DATA_COLUMN_reg_15_inst : FD1 port map( D => n7949, CP => CLK_I, Q => 
                           v_DATA_COLUMN_15_port, QN => n_3128);
   v_DATA_COLUMN_reg_16_inst : FD1 port map( D => n4331, CP => CLK_I, Q => 
                           v_DATA_COLUMN_16_port, QN => n_3129);
   v_DATA_COLUMN_reg_17_inst : FD1 port map( D => n7973, CP => CLK_I, Q => 
                           v_DATA_COLUMN_17_port, QN => n_3130);
   v_DATA_COLUMN_reg_18_inst : FD1 port map( D => n7968, CP => CLK_I, Q => 
                           v_DATA_COLUMN_18_port, QN => n_3131);
   v_DATA_COLUMN_reg_19_inst : FD1 port map( D => n7964, CP => CLK_I, Q => 
                           v_DATA_COLUMN_19_port, QN => n_3132);
   v_DATA_COLUMN_reg_20_inst : FD1 port map( D => n7960, CP => CLK_I, Q => 
                           v_DATA_COLUMN_20_port, QN => n_3133);
   v_DATA_COLUMN_reg_21_inst : FD1 port map( D => n7956, CP => CLK_I, Q => 
                           v_DATA_COLUMN_21_port, QN => n_3134);
   v_DATA_COLUMN_reg_22_inst : FD1 port map( D => n7952, CP => CLK_I, Q => 
                           v_DATA_COLUMN_22_port, QN => n_3135);
   v_DATA_COLUMN_reg_23_inst : FD1 port map( D => n7948, CP => CLK_I, Q => 
                           v_DATA_COLUMN_23_port, QN => n_3136);
   v_DATA_COLUMN_reg_0_inst : FD1 port map( D => n4323, CP => CLK_I, Q => 
                           v_DATA_COLUMN_0_port, QN => n_3137);
   v_DATA_COLUMN_reg_1_inst : FD1 port map( D => n7972, CP => CLK_I, Q => 
                           v_DATA_COLUMN_1_port, QN => n_3138);
   v_DATA_COLUMN_reg_2_inst : FD1 port map( D => n7966, CP => CLK_I, Q => 
                           v_DATA_COLUMN_2_port, QN => n_3139);
   v_DATA_COLUMN_reg_3_inst : FD1 port map( D => n7962, CP => CLK_I, Q => 
                           v_DATA_COLUMN_3_port, QN => n_3140);
   v_DATA_COLUMN_reg_4_inst : FD1 port map( D => n7958, CP => CLK_I, Q => 
                           v_DATA_COLUMN_4_port, QN => n_3141);
   v_DATA_COLUMN_reg_5_inst : FD1 port map( D => n7954, CP => CLK_I, Q => 
                           v_DATA_COLUMN_5_port, QN => n_3142);
   v_DATA_COLUMN_reg_6_inst : FD1 port map( D => n7950, CP => CLK_I, Q => 
                           v_DATA_COLUMN_6_port, QN => n_3143);
   v_DATA_COLUMN_reg_7_inst : FD1 port map( D => n7946, CP => CLK_I, Q => 
                           v_DATA_COLUMN_7_port, QN => n_3144);
   FF_VALID_DATA_reg : FD1 port map( D => n4315, CP => CLK_I, Q => n7886, QN =>
                           n4432);
   LAST_ROUND_reg : FD1 port map( D => n4314, CP => CLK_I, Q => n_3145, QN => 
                           n4400);
   v_CALCULATION_CNTR_reg_0_inst : FD1 port map( D => n4313, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_0_port, QN => n4399);
   v_CALCULATION_CNTR_reg_1_inst : FD1 port map( D => n4312, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_1_port, QN => n4405);
   v_CALCULATION_CNTR_reg_2_inst : FD1 port map( D => n4311, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_2_port, QN => n_3146);
   v_CALCULATION_CNTR_reg_3_inst : FD1 port map( D => n4310, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_3_port, QN => n4401);
   v_CALCULATION_CNTR_reg_4_inst : FD1 port map( D => n4309, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_4_port, QN => n4416);
   v_CALCULATION_CNTR_reg_5_inst : FD1 port map( D => n7977, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_5_port, QN => n_3147);
   v_CALCULATION_CNTR_reg_6_inst : FD1 port map( D => n7976, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_6_port, QN => n4417);
   v_CALCULATION_CNTR_reg_7_inst : FD1 port map( D => n7975, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_7_port, QN => n_3148);
   FF_GET_KEY_reg : FD1 port map( D => n4305, CP => CLK_I, Q => n7896, QN => 
                           n_3149);
   SRAM_WREN0_reg : FD1 port map( D => n4304, CP => CLK_I, Q => n7891, QN => 
                           n_3150);
   i_RAM_ADDR_WR0_reg_0_inst : FD1 port map( D => n4303, CP => CLK_I, Q => 
                           n7885, QN => n4433);
   i_RAM_ADDR_WR0_reg_1_inst : FD1 port map( D => n7974, CP => CLK_I, Q => 
                           n7884, QN => n4414);
   v_KEY_NUMB_reg_5_inst : FD1 port map( D => n4301, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_5_port, QN => n3947);
   v_KEY_NUMB_reg_0_inst : FD1 port map( D => n4300, CP => CLK_I, Q => 
                           v_KEY_NUMB_0_port, QN => n4419);
   v_KEY_NUMB_reg_1_inst : FD1 port map( D => n4299, CP => CLK_I, Q => 
                           v_KEY_NUMB_1_port, QN => n4435);
   v_KEY_NUMB_reg_2_inst : FD1 port map( D => n4298, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_2_port, QN => n4411);
   v_KEY_NUMB_reg_3_inst : FD1 port map( D => n4297, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_3_port, QN => n4429);
   v_KEY_NUMB_reg_4_inst : FD1 port map( D => n4296, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_4_port, QN => n_3151);
   i_RAM_ADDR_RD0_reg_0_inst : FD1 port map( D => n4295, CP => CLK_I, Q => 
                           n7888, QN => n4434);
   i_RAM_ADDR_RD0_reg_1_inst : FD1 port map( D => n4294, CP => CLK_I, Q => 
                           n7887, QN => n4415);
   CALCULATION_reg : FD1 port map( D => n4293, CP => CLK_I, Q => n7945, QN => 
                           n4431);
   i_ROUND_reg_0_inst : FD1 port map( D => n4292, CP => CLK_I, Q => n7895, QN 
                           => n4436);
   i_ROUND_reg_1_inst : FD1 port map( D => n4291, CP => CLK_I, Q => n7892, QN 
                           => n4369);
   i_ROUND_reg_2_inst : FD1 port map( D => n4290, CP => CLK_I, Q => n7893, QN 
                           => n4430);
   i_ROUND_reg_3_inst : FD1 port map( D => n4289, CP => CLK_I, Q => n7894, QN 
                           => n_3152);
   STATE_TABLE1_reg_0_7_inst : FD1 port map( D => n4288, CP => CLK_I, Q => 
                           n7851, QN => n_3153);
   STATE_TABLE1_reg_0_6_inst : FD1 port map( D => n4287, CP => CLK_I, Q => 
                           n7850, QN => n_3154);
   STATE_TABLE1_reg_0_5_inst : FD1 port map( D => n4286, CP => CLK_I, Q => 
                           n7849, QN => n_3155);
   STATE_TABLE1_reg_0_4_inst : FD1 port map( D => n4285, CP => CLK_I, Q => 
                           n7852, QN => n_3156);
   STATE_TABLE1_reg_0_3_inst : FD1 port map( D => n4284, CP => CLK_I, Q => 
                           n7859, QN => n_3157);
   STATE_TABLE1_reg_0_2_inst : FD1 port map( D => n4283, CP => CLK_I, Q => 
                           n7867, QN => n_3158);
   STATE_TABLE1_reg_0_1_inst : FD1 port map( D => n4282, CP => CLK_I, Q => 
                           n7853, QN => n_3159);
   STATE_TABLE1_reg_0_0_inst : FD1 port map( D => n4281, CP => CLK_I, Q => 
                           n7858, QN => n_3160);
   STATE_TABLE1_reg_1_7_inst : FD1 port map( D => n4280, CP => CLK_I, Q => 
                           n7848, QN => n_3161);
   STATE_TABLE1_reg_1_6_inst : FD1 port map( D => n4279, CP => CLK_I, Q => 
                           n7847, QN => n_3162);
   STATE_TABLE1_reg_1_5_inst : FD1 port map( D => n4278, CP => CLK_I, Q => 
                           n7877, QN => n_3163);
   STATE_TABLE1_reg_1_4_inst : FD1 port map( D => n4277, CP => CLK_I, Q => 
                           n7846, QN => n_3164);
   STATE_TABLE1_reg_1_3_inst : FD1 port map( D => n4276, CP => CLK_I, Q => 
                           n7845, QN => n_3165);
   STATE_TABLE1_reg_1_2_inst : FD1 port map( D => n4275, CP => CLK_I, Q => 
                           n7844, QN => n_3166);
   STATE_TABLE1_reg_1_1_inst : FD1 port map( D => n4274, CP => CLK_I, Q => 
                           n7866, QN => n_3167);
   STATE_TABLE1_reg_1_0_inst : FD1 port map( D => n4273, CP => CLK_I, Q => 
                           n7876, QN => n_3168);
   STATE_TABLE1_reg_2_7_inst : FD1 port map( D => n4272, CP => CLK_I, Q => 
                           n7897, QN => n4462);
   STATE_TABLE1_reg_2_6_inst : FD1 port map( D => n4271, CP => CLK_I, Q => 
                           n7903, QN => n4466);
   STATE_TABLE1_reg_2_5_inst : FD1 port map( D => n4270, CP => CLK_I, Q => 
                           n7909, QN => n4470);
   STATE_TABLE1_reg_2_4_inst : FD1 port map( D => n4269, CP => CLK_I, Q => 
                           n7915, QN => n4474);
   STATE_TABLE1_reg_2_3_inst : FD1 port map( D => n4268, CP => CLK_I, Q => 
                           n7921, QN => n4478);
   STATE_TABLE1_reg_2_2_inst : FD1 port map( D => n4267, CP => CLK_I, Q => 
                           n7927, QN => n4482);
   STATE_TABLE1_reg_2_1_inst : FD1 port map( D => n4266, CP => CLK_I, Q => 
                           n7933, QN => n4427);
   STATE_TABLE1_reg_2_0_inst : FD1 port map( D => n4265, CP => CLK_I, Q => 
                           n7939, QN => n4488);
   STATE_TABLE1_reg_3_7_inst : FD1 port map( D => n4264, CP => CLK_I, Q => 
                           n7898, QN => n4464);
   STATE_TABLE1_reg_3_6_inst : FD1 port map( D => n4263, CP => CLK_I, Q => 
                           n7904, QN => n4468);
   STATE_TABLE1_reg_3_5_inst : FD1 port map( D => n4262, CP => CLK_I, Q => 
                           n7910, QN => n4472);
   STATE_TABLE1_reg_3_4_inst : FD1 port map( D => n4261, CP => CLK_I, Q => 
                           n7916, QN => n4476);
   STATE_TABLE1_reg_3_3_inst : FD1 port map( D => n4260, CP => CLK_I, Q => 
                           n7922, QN => n4480);
   STATE_TABLE1_reg_3_2_inst : FD1 port map( D => n4259, CP => CLK_I, Q => 
                           n7928, QN => n4484);
   STATE_TABLE1_reg_3_1_inst : FD1 port map( D => n4258, CP => CLK_I, Q => 
                           n7934, QN => n4428);
   STATE_TABLE1_reg_3_0_inst : FD1 port map( D => n4257, CP => CLK_I, Q => 
                           n7940, QN => n4490);
   STATE_TABLE1_reg_4_7_inst : FD1 port map( D => n4256, CP => CLK_I, Q => 
                           n7899, QN => n4384);
   STATE_TABLE1_reg_4_6_inst : FD1 port map( D => n4255, CP => CLK_I, Q => 
                           n7905, QN => n4386);
   STATE_TABLE1_reg_4_5_inst : FD1 port map( D => n4254, CP => CLK_I, Q => 
                           n7911, QN => n4378);
   STATE_TABLE1_reg_4_4_inst : FD1 port map( D => n4253, CP => CLK_I, Q => 
                           n7917, QN => n4388);
   STATE_TABLE1_reg_4_3_inst : FD1 port map( D => n4252, CP => CLK_I, Q => 
                           n7923, QN => n4380);
   STATE_TABLE1_reg_4_2_inst : FD1 port map( D => n4251, CP => CLK_I, Q => 
                           n7929, QN => n4382);
   STATE_TABLE1_reg_4_1_inst : FD1 port map( D => n4250, CP => CLK_I, Q => 
                           n7935, QN => n4391);
   STATE_TABLE1_reg_4_0_inst : FD1 port map( D => n4249, CP => CLK_I, Q => 
                           n7941, QN => n4392);
   STATE_TABLE1_reg_5_7_inst : FD1 port map( D => n4248, CP => CLK_I, Q => 
                           n7843, QN => n_3169);
   STATE_TABLE1_reg_5_6_inst : FD1 port map( D => n4247, CP => CLK_I, Q => 
                           n7842, QN => n_3170);
   STATE_TABLE1_reg_5_5_inst : FD1 port map( D => n4246, CP => CLK_I, Q => 
                           n7880, QN => n_3171);
   STATE_TABLE1_reg_5_4_inst : FD1 port map( D => n4245, CP => CLK_I, Q => 
                           n7841, QN => n_3172);
   STATE_TABLE1_reg_5_3_inst : FD1 port map( D => n4244, CP => CLK_I, Q => 
                           n7840, QN => n_3173);
   STATE_TABLE1_reg_5_2_inst : FD1 port map( D => n4243, CP => CLK_I, Q => 
                           n7839, QN => n_3174);
   STATE_TABLE1_reg_5_1_inst : FD1 port map( D => n4242, CP => CLK_I, Q => 
                           n7838, QN => n_3175);
   STATE_TABLE1_reg_5_0_inst : FD1 port map( D => n4241, CP => CLK_I, Q => 
                           n7879, QN => n_3176);
   STATE_TABLE1_reg_6_7_inst : FD1 port map( D => n4240, CP => CLK_I, Q => 
                           n7837, QN => n_3177);
   STATE_TABLE1_reg_6_6_inst : FD1 port map( D => n4239, CP => CLK_I, Q => 
                           n7836, QN => n_3178);
   STATE_TABLE1_reg_6_5_inst : FD1 port map( D => n4238, CP => CLK_I, Q => 
                           n7835, QN => n_3179);
   STATE_TABLE1_reg_6_4_inst : FD1 port map( D => n4237, CP => CLK_I, Q => 
                           n7834, QN => n_3180);
   STATE_TABLE1_reg_6_3_inst : FD1 port map( D => n4236, CP => CLK_I, Q => 
                           n7864, QN => n_3181);
   STATE_TABLE1_reg_6_2_inst : FD1 port map( D => n4235, CP => CLK_I, Q => 
                           n7872, QN => n_3182);
   STATE_TABLE1_reg_6_1_inst : FD1 port map( D => n4234, CP => CLK_I, Q => 
                           n7833, QN => n_3183);
   STATE_TABLE1_reg_6_0_inst : FD1 port map( D => n4233, CP => CLK_I, Q => 
                           n7878, QN => n_3184);
   STATE_TABLE1_reg_7_7_inst : FD1 port map( D => n4232, CP => CLK_I, Q => 
                           n7832, QN => n4463);
   STATE_TABLE1_reg_7_6_inst : FD1 port map( D => n4231, CP => CLK_I, Q => 
                           n7831, QN => n4467);
   STATE_TABLE1_reg_7_5_inst : FD1 port map( D => n4230, CP => CLK_I, Q => 
                           n7830, QN => n4471);
   STATE_TABLE1_reg_7_4_inst : FD1 port map( D => n4229, CP => CLK_I, Q => 
                           n7857, QN => n4475);
   STATE_TABLE1_reg_7_3_inst : FD1 port map( D => n4228, CP => CLK_I, Q => 
                           n7829, QN => n4479);
   STATE_TABLE1_reg_7_2_inst : FD1 port map( D => n4227, CP => CLK_I, Q => 
                           n7871, QN => n4483);
   STATE_TABLE1_reg_7_1_inst : FD1 port map( D => n4226, CP => CLK_I, Q => 
                           n7863, QN => n4486);
   STATE_TABLE1_reg_7_0_inst : FD1 port map( D => n4225, CP => CLK_I, Q => 
                           n7828, QN => n4489);
   STATE_TABLE1_reg_8_7_inst : FD1 port map( D => n4224, CP => CLK_I, Q => 
                           n7827, QN => n_3185);
   STATE_TABLE1_reg_8_6_inst : FD1 port map( D => n4223, CP => CLK_I, Q => 
                           n7826, QN => n_3186);
   STATE_TABLE1_reg_8_5_inst : FD1 port map( D => n4222, CP => CLK_I, Q => 
                           n7825, QN => n_3187);
   STATE_TABLE1_reg_8_4_inst : FD1 port map( D => n4221, CP => CLK_I, Q => 
                           n7854, QN => n_3188);
   STATE_TABLE1_reg_8_3_inst : FD1 port map( D => n4220, CP => CLK_I, Q => 
                           n7862, QN => n_3189);
   STATE_TABLE1_reg_8_2_inst : FD1 port map( D => n4219, CP => CLK_I, Q => 
                           n7870, QN => n_3190);
   STATE_TABLE1_reg_8_1_inst : FD1 port map( D => n4218, CP => CLK_I, Q => 
                           n7855, QN => n_3191);
   STATE_TABLE1_reg_8_0_inst : FD1 port map( D => n4217, CP => CLK_I, Q => 
                           n7861, QN => n_3192);
   STATE_TABLE1_reg_9_7_inst : FD1 port map( D => n4216, CP => CLK_I, Q => 
                           n7824, QN => n_3193);
   STATE_TABLE1_reg_9_6_inst : FD1 port map( D => n4215, CP => CLK_I, Q => 
                           n7823, QN => n_3194);
   STATE_TABLE1_reg_9_5_inst : FD1 port map( D => n4214, CP => CLK_I, Q => 
                           n7882, QN => n_3195);
   STATE_TABLE1_reg_9_4_inst : FD1 port map( D => n4213, CP => CLK_I, Q => 
                           n7822, QN => n_3196);
   STATE_TABLE1_reg_9_3_inst : FD1 port map( D => n4212, CP => CLK_I, Q => 
                           n7821, QN => n_3197);
   STATE_TABLE1_reg_9_2_inst : FD1 port map( D => n4211, CP => CLK_I, Q => 
                           n7820, QN => n_3198);
   STATE_TABLE1_reg_9_1_inst : FD1 port map( D => n4210, CP => CLK_I, Q => 
                           n7868, QN => n_3199);
   STATE_TABLE1_reg_9_0_inst : FD1 port map( D => n4209, CP => CLK_I, Q => 
                           n7881, QN => n_3200);
   STATE_TABLE1_reg_10_7_inst : FD1 port map( D => n4208, CP => CLK_I, Q => 
                           n7901, QN => n4465);
   STATE_TABLE1_reg_10_6_inst : FD1 port map( D => n4207, CP => CLK_I, Q => 
                           n7907, QN => n4469);
   STATE_TABLE1_reg_10_5_inst : FD1 port map( D => n4206, CP => CLK_I, Q => 
                           n7913, QN => n4473);
   STATE_TABLE1_reg_10_4_inst : FD1 port map( D => n4205, CP => CLK_I, Q => 
                           n7919, QN => n4477);
   STATE_TABLE1_reg_10_3_inst : FD1 port map( D => n4204, CP => CLK_I, Q => 
                           n7925, QN => n4481);
   STATE_TABLE1_reg_10_2_inst : FD1 port map( D => n4203, CP => CLK_I, Q => 
                           n7931, QN => n4485);
   STATE_TABLE1_reg_10_1_inst : FD1 port map( D => n4202, CP => CLK_I, Q => 
                           n7937, QN => n4487);
   STATE_TABLE1_reg_10_0_inst : FD1 port map( D => n4201, CP => CLK_I, Q => 
                           n7943, QN => n4491);
   STATE_TABLE1_reg_11_7_inst : FD1 port map( D => n4200, CP => CLK_I, Q => 
                           n7819, QN => n_3201);
   STATE_TABLE1_reg_11_6_inst : FD1 port map( D => n4199, CP => CLK_I, Q => 
                           n7818, QN => n_3202);
   STATE_TABLE1_reg_11_5_inst : FD1 port map( D => n4198, CP => CLK_I, Q => 
                           n7817, QN => n_3203);
   STATE_TABLE1_reg_11_4_inst : FD1 port map( D => n4197, CP => CLK_I, Q => 
                           n7856, QN => n_3204);
   STATE_TABLE1_reg_11_3_inst : FD1 port map( D => n4196, CP => CLK_I, Q => 
                           n7816, QN => n_3205);
   STATE_TABLE1_reg_11_2_inst : FD1 port map( D => n4195, CP => CLK_I, Q => 
                           n7869, QN => n_3206);
   STATE_TABLE1_reg_11_1_inst : FD1 port map( D => n4194, CP => CLK_I, Q => 
                           n7860, QN => n_3207);
   STATE_TABLE1_reg_11_0_inst : FD1 port map( D => n4193, CP => CLK_I, Q => 
                           n7815, QN => n_3208);
   STATE_TABLE1_reg_12_7_inst : FD1 port map( D => n4192, CP => CLK_I, Q => 
                           n7902, QN => n4385);
   STATE_TABLE1_reg_12_6_inst : FD1 port map( D => n4191, CP => CLK_I, Q => 
                           n7908, QN => n4387);
   STATE_TABLE1_reg_12_5_inst : FD1 port map( D => n4190, CP => CLK_I, Q => 
                           n7914, QN => n4379);
   STATE_TABLE1_reg_12_4_inst : FD1 port map( D => n4189, CP => CLK_I, Q => 
                           n7920, QN => n4389);
   STATE_TABLE1_reg_12_3_inst : FD1 port map( D => n4188, CP => CLK_I, Q => 
                           n7926, QN => n4381);
   STATE_TABLE1_reg_12_2_inst : FD1 port map( D => n4187, CP => CLK_I, Q => 
                           n7932, QN => n4390);
   STATE_TABLE1_reg_12_1_inst : FD1 port map( D => n4186, CP => CLK_I, Q => 
                           n7938, QN => n4383);
   STATE_TABLE1_reg_12_0_inst : FD1 port map( D => n4185, CP => CLK_I, Q => 
                           n7944, QN => n4393);
   STATE_TABLE1_reg_13_7_inst : FD1 port map( D => n4184, CP => CLK_I, Q => 
                           n7814, QN => n_3209);
   STATE_TABLE1_reg_13_6_inst : FD1 port map( D => n4183, CP => CLK_I, Q => 
                           n7813, QN => n_3210);
   STATE_TABLE1_reg_13_5_inst : FD1 port map( D => n4182, CP => CLK_I, Q => 
                           n7883, QN => n_3211);
   STATE_TABLE1_reg_13_4_inst : FD1 port map( D => n4181, CP => CLK_I, Q => 
                           n7812, QN => n_3212);
   STATE_TABLE1_reg_13_3_inst : FD1 port map( D => n4180, CP => CLK_I, Q => 
                           n7811, QN => n_3213);
   STATE_TABLE1_reg_13_2_inst : FD1 port map( D => n4179, CP => CLK_I, Q => 
                           n7810, QN => n_3214);
   STATE_TABLE1_reg_13_1_inst : FD1 port map( D => n4178, CP => CLK_I, Q => 
                           n7809, QN => n_3215);
   STATE_TABLE1_reg_13_0_inst : FD1 port map( D => n4177, CP => CLK_I, Q => 
                           n7808, QN => n_3216);
   STATE_TABLE1_reg_14_7_inst : FD1 port map( D => n4176, CP => CLK_I, Q => 
                           n7875, QN => n_3217);
   STATE_TABLE1_reg_14_6_inst : FD1 port map( D => n4175, CP => CLK_I, Q => 
                           n7889, QN => n_3218);
   STATE_TABLE1_reg_14_5_inst : FD1 port map( D => n4174, CP => CLK_I, Q => 
                           n7890, QN => n_3219);
   STATE_TABLE1_reg_14_4_inst : FD1 port map( D => n4173, CP => CLK_I, Q => 
                           n7807, QN => n_3220);
   STATE_TABLE1_reg_14_3_inst : FD1 port map( D => n4172, CP => CLK_I, Q => 
                           n7865, QN => n_3221);
   STATE_TABLE1_reg_14_2_inst : FD1 port map( D => n4171, CP => CLK_I, Q => 
                           n7874, QN => n_3222);
   STATE_TABLE1_reg_14_1_inst : FD1 port map( D => n4170, CP => CLK_I, Q => 
                           n7873, QN => n_3223);
   STATE_TABLE1_reg_14_0_inst : FD1 port map( D => n4169, CP => CLK_I, Q => 
                           n7806, QN => n_3224);
   STATE_TABLE1_reg_15_7_inst : FD1 port map( D => n4168, CP => CLK_I, Q => 
                           n7900, QN => n_3225);
   STATE_TABLE1_reg_15_6_inst : FD1 port map( D => n4167, CP => CLK_I, Q => 
                           n7906, QN => n_3226);
   STATE_TABLE1_reg_15_5_inst : FD1 port map( D => n4166, CP => CLK_I, Q => 
                           n7912, QN => n_3227);
   v_RAM_IN0_reg_24_inst : FD1 port map( D => n4165, CP => CLK_I, Q => 
                           v_RAM_IN0_24_port, QN => n4371);
   t_STATE_RAM0_reg_0_24_inst : FD1 port map( D => n4164, CP => CLK_I, Q => 
                           n_3228, QN => n4420);
   t_STATE_RAM0_reg_1_24_inst : FD1 port map( D => n4163, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_24_port, QN => n_3229);
   t_STATE_RAM0_reg_2_24_inst : FD1 port map( D => n4162, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_24_port, QN => n_3230);
   t_STATE_RAM0_reg_3_24_inst : FD1 port map( D => n4161, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_24_port, QN => n_3231);
   v_RAM_OUT0_reg_24_inst : FD1 port map( D => n4160, CP => CLK_I, Q => 
                           v_RAM_OUT0_24_port, QN => n4355);
   STATE_TABLE1_reg_15_4_inst : FD1 port map( D => n4159, CP => CLK_I, Q => 
                           n7918, QN => n_3232);
   v_RAM_IN0_reg_31_inst : FD1 port map( D => n4158, CP => CLK_I, Q => 
                           v_RAM_IN0_31_port, QN => n_3233);
   t_STATE_RAM0_reg_0_31_inst : FD1 port map( D => n4157, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_31_port, QN => n4437);
   t_STATE_RAM0_reg_1_31_inst : FD1 port map( D => n4156, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_31_port, QN => n_3234);
   t_STATE_RAM0_reg_2_31_inst : FD1 port map( D => n4155, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_31_port, QN => n_3235);
   t_STATE_RAM0_reg_3_31_inst : FD1 port map( D => n4154, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_31_port, QN => n_3236);
   v_RAM_OUT0_reg_31_inst : FD1 port map( D => n4153, CP => CLK_I, Q => 
                           v_RAM_OUT0_31_port, QN => n4396);
   v_RAM_IN0_reg_23_inst : FD1 port map( D => n4152, CP => CLK_I, Q => 
                           v_RAM_IN0_23_port, QN => n4372);
   t_STATE_RAM0_reg_0_23_inst : FD1 port map( D => n4151, CP => CLK_I, Q => 
                           n_3237, QN => n4421);
   t_STATE_RAM0_reg_1_23_inst : FD1 port map( D => n4150, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_23_port, QN => n_3238);
   t_STATE_RAM0_reg_2_23_inst : FD1 port map( D => n4149, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_23_port, QN => n_3239);
   t_STATE_RAM0_reg_3_23_inst : FD1 port map( D => n4148, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_23_port, QN => n_3240);
   v_RAM_OUT0_reg_23_inst : FD1 port map( D => n4147, CP => CLK_I, Q => 
                           v_RAM_OUT0_23_port, QN => n4395);
   v_RAM_IN0_reg_15_inst : FD1 port map( D => n4146, CP => CLK_I, Q => 
                           v_RAM_IN0_15_port, QN => n_3241);
   t_STATE_RAM0_reg_0_15_inst : FD1 port map( D => n4145, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_15_port, QN => n4438);
   t_STATE_RAM0_reg_1_15_inst : FD1 port map( D => n4144, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_15_port, QN => n_3242);
   t_STATE_RAM0_reg_2_15_inst : FD1 port map( D => n4143, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_15_port, QN => n_3243);
   t_STATE_RAM0_reg_3_15_inst : FD1 port map( D => n4142, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_15_port, QN => n_3244);
   v_RAM_OUT0_reg_15_inst : FD1 port map( D => n4141, CP => CLK_I, Q => 
                           v_RAM_OUT0_15_port, QN => n4397);
   v_RAM_IN0_reg_7_inst : FD1 port map( D => n4140, CP => CLK_I, Q => 
                           v_RAM_IN0_7_port, QN => n_3245);
   t_STATE_RAM0_reg_0_7_inst : FD1 port map( D => n4139, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_7_port, QN => n4439);
   t_STATE_RAM0_reg_1_7_inst : FD1 port map( D => n4138, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_7_port, QN => n_3246);
   t_STATE_RAM0_reg_2_7_inst : FD1 port map( D => n4137, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_7_port, QN => n_3247);
   t_STATE_RAM0_reg_3_7_inst : FD1 port map( D => n4136, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_7_port, QN => n_3248);
   v_RAM_OUT0_reg_7_inst : FD1 port map( D => n4135, CP => CLK_I, Q => 
                           v_RAM_OUT0_7_port, QN => n4394);
   STATE_TABLE1_reg_15_3_inst : FD1 port map( D => n4134, CP => CLK_I, Q => 
                           n7924, QN => n_3249);
   v_RAM_IN0_reg_30_inst : FD1 port map( D => n4133, CP => CLK_I, Q => 
                           v_RAM_IN0_30_port, QN => n4373);
   t_STATE_RAM0_reg_0_30_inst : FD1 port map( D => n4132, CP => CLK_I, Q => 
                           n_3250, QN => n4422);
   t_STATE_RAM0_reg_1_30_inst : FD1 port map( D => n4131, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_30_port, QN => n_3251);
   t_STATE_RAM0_reg_2_30_inst : FD1 port map( D => n4130, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_30_port, QN => n_3252);
   t_STATE_RAM0_reg_3_30_inst : FD1 port map( D => n4129, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_30_port, QN => n_3253);
   v_RAM_OUT0_reg_30_inst : FD1 port map( D => n4128, CP => CLK_I, Q => 
                           v_RAM_OUT0_30_port, QN => n4413);
   v_RAM_IN0_reg_22_inst : FD1 port map( D => n4127, CP => CLK_I, Q => 
                           v_RAM_IN0_22_port, QN => n4374);
   t_STATE_RAM0_reg_0_22_inst : FD1 port map( D => n4126, CP => CLK_I, Q => 
                           n_3254, QN => n4423);
   t_STATE_RAM0_reg_1_22_inst : FD1 port map( D => n4125, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_22_port, QN => n_3255);
   t_STATE_RAM0_reg_2_22_inst : FD1 port map( D => n4124, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_22_port, QN => n_3256);
   t_STATE_RAM0_reg_3_22_inst : FD1 port map( D => n4123, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_22_port, QN => n_3257);
   v_RAM_OUT0_reg_22_inst : FD1 port map( D => n4122, CP => CLK_I, Q => 
                           v_RAM_OUT0_22_port, QN => n4412);
   v_RAM_IN0_reg_14_inst : FD1 port map( D => n4121, CP => CLK_I, Q => 
                           v_RAM_IN0_14_port, QN => n4375);
   t_STATE_RAM0_reg_0_14_inst : FD1 port map( D => n4120, CP => CLK_I, Q => 
                           n_3258, QN => n4424);
   t_STATE_RAM0_reg_1_14_inst : FD1 port map( D => n4119, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_14_port, QN => n_3259);
   t_STATE_RAM0_reg_2_14_inst : FD1 port map( D => n4118, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_14_port, QN => n_3260);
   t_STATE_RAM0_reg_3_14_inst : FD1 port map( D => n4117, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_14_port, QN => n_3261);
   v_RAM_OUT0_reg_14_inst : FD1 port map( D => n4116, CP => CLK_I, Q => 
                           v_RAM_OUT0_14_port, QN => n4366);
   v_RAM_IN0_reg_6_inst : FD1 port map( D => n4115, CP => CLK_I, Q => 
                           v_RAM_IN0_6_port, QN => n4376);
   t_STATE_RAM0_reg_0_6_inst : FD1 port map( D => n4114, CP => CLK_I, Q => 
                           n_3262, QN => n4425);
   t_STATE_RAM0_reg_1_6_inst : FD1 port map( D => n4113, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_6_port, QN => n_3263);
   t_STATE_RAM0_reg_2_6_inst : FD1 port map( D => n4112, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_6_port, QN => n_3264);
   t_STATE_RAM0_reg_3_6_inst : FD1 port map( D => n4111, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_6_port, QN => n_3265);
   v_RAM_OUT0_reg_6_inst : FD1 port map( D => n4110, CP => CLK_I, Q => 
                           v_RAM_OUT0_6_port, QN => n4407);
   STATE_TABLE1_reg_15_2_inst : FD1 port map( D => n4109, CP => CLK_I, Q => 
                           n7930, QN => n_3266);
   v_RAM_IN0_reg_21_inst : FD1 port map( D => n4108, CP => CLK_I, Q => 
                           v_RAM_IN0_21_port, QN => n_3267);
   t_STATE_RAM0_reg_0_21_inst : FD1 port map( D => n4107, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_21_port, QN => n4440);
   t_STATE_RAM0_reg_1_21_inst : FD1 port map( D => n4106, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_21_port, QN => n_3268);
   t_STATE_RAM0_reg_2_21_inst : FD1 port map( D => n4105, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_21_port, QN => n_3269);
   t_STATE_RAM0_reg_3_21_inst : FD1 port map( D => n4104, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_21_port, QN => n_3270);
   v_RAM_OUT0_reg_21_inst : FD1 port map( D => n4103, CP => CLK_I, Q => 
                           v_RAM_OUT0_21_port, QN => n4403);
   v_RAM_IN0_reg_13_inst : FD1 port map( D => n4102, CP => CLK_I, Q => 
                           v_RAM_IN0_13_port, QN => n_3271);
   t_STATE_RAM0_reg_0_13_inst : FD1 port map( D => n4101, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_13_port, QN => n4441);
   t_STATE_RAM0_reg_1_13_inst : FD1 port map( D => n4100, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_13_port, QN => n_3272);
   t_STATE_RAM0_reg_2_13_inst : FD1 port map( D => n4099, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_13_port, QN => n_3273);
   t_STATE_RAM0_reg_3_13_inst : FD1 port map( D => n4098, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_13_port, QN => n_3274);
   v_RAM_OUT0_reg_13_inst : FD1 port map( D => n4097, CP => CLK_I, Q => 
                           v_RAM_OUT0_13_port, QN => n4353);
   v_RAM_IN0_reg_29_inst : FD1 port map( D => n4096, CP => CLK_I, Q => 
                           v_RAM_IN0_29_port, QN => n_3275);
   t_STATE_RAM0_reg_0_29_inst : FD1 port map( D => n4095, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_29_port, QN => n4442);
   t_STATE_RAM0_reg_1_29_inst : FD1 port map( D => n4094, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_29_port, QN => n_3276);
   t_STATE_RAM0_reg_2_29_inst : FD1 port map( D => n4093, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_29_port, QN => n_3277);
   t_STATE_RAM0_reg_3_29_inst : FD1 port map( D => n4092, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_29_port, QN => n_3278);
   v_RAM_OUT0_reg_29_inst : FD1 port map( D => n4091, CP => CLK_I, Q => 
                           v_RAM_OUT0_29_port, QN => n4404);
   v_RAM_IN0_reg_5_inst : FD1 port map( D => n4090, CP => CLK_I, Q => 
                           v_RAM_IN0_5_port, QN => n_3279);
   t_STATE_RAM0_reg_0_5_inst : FD1 port map( D => n4089, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_5_port, QN => n4443);
   t_STATE_RAM0_reg_1_5_inst : FD1 port map( D => n4088, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_5_port, QN => n_3280);
   t_STATE_RAM0_reg_2_5_inst : FD1 port map( D => n4087, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_5_port, QN => n_3281);
   t_STATE_RAM0_reg_3_5_inst : FD1 port map( D => n4086, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_5_port, QN => n_3282);
   v_RAM_OUT0_reg_5_inst : FD1 port map( D => n4085, CP => CLK_I, Q => 
                           v_RAM_OUT0_5_port, QN => n4402);
   v_RAM_IN0_reg_2_inst : FD1 port map( D => n4084, CP => CLK_I, Q => 
                           v_RAM_IN0_2_port, QN => n_3283);
   t_STATE_RAM0_reg_0_2_inst : FD1 port map( D => n4083, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_2_port, QN => n4444);
   t_STATE_RAM0_reg_1_2_inst : FD1 port map( D => n4082, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_2_port, QN => n_3284);
   t_STATE_RAM0_reg_2_2_inst : FD1 port map( D => n4081, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_2_port, QN => n_3285);
   t_STATE_RAM0_reg_3_2_inst : FD1 port map( D => n4080, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_2_port, QN => n_3286);
   v_RAM_OUT0_reg_2_inst : FD1 port map( D => n4079, CP => CLK_I, Q => 
                           v_RAM_OUT0_2_port, QN => n4360);
   STATE_TABLE1_reg_15_1_inst : FD1 port map( D => n4078, CP => CLK_I, Q => 
                           n7936, QN => n_3287);
   v_RAM_IN0_reg_18_inst : FD1 port map( D => n4077, CP => CLK_I, Q => 
                           v_RAM_IN0_18_port, QN => n_3288);
   t_STATE_RAM0_reg_0_18_inst : FD1 port map( D => n4076, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_18_port, QN => n4445);
   t_STATE_RAM0_reg_1_18_inst : FD1 port map( D => n4075, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_18_port, QN => n_3289);
   t_STATE_RAM0_reg_2_18_inst : FD1 port map( D => n4074, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_18_port, QN => n_3290);
   t_STATE_RAM0_reg_3_18_inst : FD1 port map( D => n4073, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_18_port, QN => n_3291);
   v_RAM_OUT0_reg_18_inst : FD1 port map( D => n4072, CP => CLK_I, Q => 
                           v_RAM_OUT0_18_port, QN => n4358);
   v_RAM_IN0_reg_9_inst : FD1 port map( D => n4071, CP => CLK_I, Q => 
                           v_RAM_IN0_9_port, QN => n_3292);
   t_STATE_RAM0_reg_0_9_inst : FD1 port map( D => n4070, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_9_port, QN => n4446);
   t_STATE_RAM0_reg_1_9_inst : FD1 port map( D => n4069, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_9_port, QN => n_3293);
   t_STATE_RAM0_reg_2_9_inst : FD1 port map( D => n4068, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_9_port, QN => n_3294);
   t_STATE_RAM0_reg_3_9_inst : FD1 port map( D => n4067, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_9_port, QN => n_3295);
   v_RAM_OUT0_reg_9_inst : FD1 port map( D => n4066, CP => CLK_I, Q => 
                           v_RAM_OUT0_9_port, QN => n4361);
   v_RAM_IN0_reg_28_inst : FD1 port map( D => n4065, CP => CLK_I, Q => 
                           v_RAM_IN0_28_port, QN => n_3296);
   t_STATE_RAM0_reg_0_28_inst : FD1 port map( D => n4064, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_28_port, QN => n4447);
   t_STATE_RAM0_reg_1_28_inst : FD1 port map( D => n4063, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_28_port, QN => n_3297);
   t_STATE_RAM0_reg_2_28_inst : FD1 port map( D => n4062, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_28_port, QN => n_3298);
   t_STATE_RAM0_reg_3_28_inst : FD1 port map( D => n4061, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_28_port, QN => n_3299);
   v_RAM_OUT0_reg_28_inst : FD1 port map( D => n4060, CP => CLK_I, Q => 
                           v_RAM_OUT0_28_port, QN => n4410);
   v_RAM_IN0_reg_12_inst : FD1 port map( D => n4059, CP => CLK_I, Q => 
                           v_RAM_IN0_12_port, QN => n_3300);
   t_STATE_RAM0_reg_0_12_inst : FD1 port map( D => n4058, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_12_port, QN => n4448);
   t_STATE_RAM0_reg_1_12_inst : FD1 port map( D => n4057, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_12_port, QN => n_3301);
   t_STATE_RAM0_reg_2_12_inst : FD1 port map( D => n4056, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_12_port, QN => n_3302);
   t_STATE_RAM0_reg_3_12_inst : FD1 port map( D => n4055, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_12_port, QN => n_3303);
   v_RAM_OUT0_reg_12_inst : FD1 port map( D => n4054, CP => CLK_I, Q => 
                           v_RAM_OUT0_12_port, QN => n4398);
   v_RAM_IN0_reg_20_inst : FD1 port map( D => n4053, CP => CLK_I, Q => 
                           v_RAM_IN0_20_port, QN => n_3304);
   t_STATE_RAM0_reg_0_20_inst : FD1 port map( D => n4052, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_20_port, QN => n4449);
   t_STATE_RAM0_reg_1_20_inst : FD1 port map( D => n4051, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_20_port, QN => n_3305);
   t_STATE_RAM0_reg_2_20_inst : FD1 port map( D => n4050, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_20_port, QN => n_3306);
   t_STATE_RAM0_reg_3_20_inst : FD1 port map( D => n4049, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_20_port, QN => n_3307);
   v_RAM_OUT0_reg_20_inst : FD1 port map( D => n4048, CP => CLK_I, Q => 
                           v_RAM_OUT0_20_port, QN => n4409);
   v_RAM_IN0_reg_4_inst : FD1 port map( D => n4047, CP => CLK_I, Q => 
                           v_RAM_IN0_4_port, QN => n_3308);
   t_STATE_RAM0_reg_0_4_inst : FD1 port map( D => n4046, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_4_port, QN => n4450);
   t_STATE_RAM0_reg_1_4_inst : FD1 port map( D => n4045, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_4_port, QN => n_3309);
   t_STATE_RAM0_reg_2_4_inst : FD1 port map( D => n4044, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_4_port, QN => n_3310);
   t_STATE_RAM0_reg_3_4_inst : FD1 port map( D => n4043, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_4_port, QN => n_3311);
   v_RAM_OUT0_reg_4_inst : FD1 port map( D => n4042, CP => CLK_I, Q => 
                           v_RAM_OUT0_4_port, QN => n4406);
   v_RAM_IN0_reg_1_inst : FD1 port map( D => n4041, CP => CLK_I, Q => 
                           v_RAM_IN0_1_port, QN => n_3312);
   t_STATE_RAM0_reg_0_1_inst : FD1 port map( D => n4040, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_1_port, QN => n4451);
   t_STATE_RAM0_reg_1_1_inst : FD1 port map( D => n4039, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_1_port, QN => n_3313);
   t_STATE_RAM0_reg_2_1_inst : FD1 port map( D => n4038, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_1_port, QN => n_3314);
   t_STATE_RAM0_reg_3_1_inst : FD1 port map( D => n4037, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_1_port, QN => n_3315);
   v_RAM_OUT0_reg_1_inst : FD1 port map( D => n4036, CP => CLK_I, Q => 
                           v_RAM_OUT0_1_port, QN => n4362);
   STATE_TABLE1_reg_15_0_inst : FD1 port map( D => n4035, CP => CLK_I, Q => 
                           n7942, QN => n_3316);
   v_RAM_IN0_reg_25_inst : FD1 port map( D => n4034, CP => CLK_I, Q => 
                           v_RAM_IN0_25_port, QN => n_3317);
   t_STATE_RAM0_reg_0_25_inst : FD1 port map( D => n4033, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_25_port, QN => n4452);
   t_STATE_RAM0_reg_1_25_inst : FD1 port map( D => n4032, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_25_port, QN => n_3318);
   t_STATE_RAM0_reg_2_25_inst : FD1 port map( D => n4031, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_25_port, QN => n_3319);
   t_STATE_RAM0_reg_3_25_inst : FD1 port map( D => n4030, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_25_port, QN => n_3320);
   v_RAM_OUT0_reg_25_inst : FD1 port map( D => n4029, CP => CLK_I, Q => 
                           v_RAM_OUT0_25_port, QN => n4364);
   v_RAM_IN0_reg_17_inst : FD1 port map( D => n4028, CP => CLK_I, Q => 
                           v_RAM_IN0_17_port, QN => n_3321);
   t_STATE_RAM0_reg_0_17_inst : FD1 port map( D => n4027, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_17_port, QN => n4453);
   t_STATE_RAM0_reg_1_17_inst : FD1 port map( D => n4026, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_17_port, QN => n_3322);
   t_STATE_RAM0_reg_2_17_inst : FD1 port map( D => n4025, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_17_port, QN => n_3323);
   t_STATE_RAM0_reg_3_17_inst : FD1 port map( D => n4024, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_17_port, QN => n_3324);
   v_RAM_OUT0_reg_17_inst : FD1 port map( D => n4023, CP => CLK_I, Q => 
                           v_RAM_OUT0_17_port, QN => n4363);
   v_RAM_IN0_reg_26_inst : FD1 port map( D => n4022, CP => CLK_I, Q => 
                           v_RAM_IN0_26_port, QN => n_3325);
   t_STATE_RAM0_reg_0_26_inst : FD1 port map( D => n4021, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_26_port, QN => n4454);
   t_STATE_RAM0_reg_1_26_inst : FD1 port map( D => n4020, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_26_port, QN => n_3326);
   t_STATE_RAM0_reg_2_26_inst : FD1 port map( D => n4019, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_26_port, QN => n_3327);
   t_STATE_RAM0_reg_3_26_inst : FD1 port map( D => n4018, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_26_port, QN => n_3328);
   v_RAM_OUT0_reg_26_inst : FD1 port map( D => n4017, CP => CLK_I, Q => 
                           v_RAM_OUT0_26_port, QN => n4359);
   v_RAM_IN0_reg_10_inst : FD1 port map( D => n4016, CP => CLK_I, Q => 
                           v_RAM_IN0_10_port, QN => n_3329);
   t_STATE_RAM0_reg_0_10_inst : FD1 port map( D => n4015, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_10_port, QN => n4455);
   t_STATE_RAM0_reg_1_10_inst : FD1 port map( D => n4014, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_10_port, QN => n_3330);
   t_STATE_RAM0_reg_2_10_inst : FD1 port map( D => n4013, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_10_port, QN => n_3331);
   t_STATE_RAM0_reg_3_10_inst : FD1 port map( D => n4012, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_10_port, QN => n_3332);
   v_RAM_OUT0_reg_10_inst : FD1 port map( D => n4011, CP => CLK_I, Q => 
                           v_RAM_OUT0_10_port, QN => n4357);
   v_RAM_IN0_reg_27_inst : FD1 port map( D => n4010, CP => CLK_I, Q => 
                           v_RAM_IN0_27_port, QN => n_3333);
   t_STATE_RAM0_reg_0_27_inst : FD1 port map( D => n4009, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_27_port, QN => n4456);
   t_STATE_RAM0_reg_1_27_inst : FD1 port map( D => n4008, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_27_port, QN => n_3334);
   t_STATE_RAM0_reg_2_27_inst : FD1 port map( D => n4007, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_27_port, QN => n_3335);
   t_STATE_RAM0_reg_3_27_inst : FD1 port map( D => n4006, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_27_port, QN => n_3336);
   v_RAM_OUT0_reg_27_inst : FD1 port map( D => n4005, CP => CLK_I, Q => 
                           v_RAM_OUT0_27_port, QN => n4368);
   v_RAM_IN0_reg_19_inst : FD1 port map( D => n4004, CP => CLK_I, Q => 
                           v_RAM_IN0_19_port, QN => n_3337);
   t_STATE_RAM0_reg_0_19_inst : FD1 port map( D => n4003, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_19_port, QN => n4457);
   t_STATE_RAM0_reg_1_19_inst : FD1 port map( D => n4002, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_19_port, QN => n_3338);
   t_STATE_RAM0_reg_2_19_inst : FD1 port map( D => n4001, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_19_port, QN => n_3339);
   t_STATE_RAM0_reg_3_19_inst : FD1 port map( D => n4000, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_19_port, QN => n_3340);
   v_RAM_OUT0_reg_19_inst : FD1 port map( D => n3999, CP => CLK_I, Q => 
                           v_RAM_OUT0_19_port, QN => n4367);
   v_RAM_IN0_reg_11_inst : FD1 port map( D => n3998, CP => CLK_I, Q => 
                           v_RAM_IN0_11_port, QN => n_3341);
   t_STATE_RAM0_reg_0_11_inst : FD1 port map( D => n3997, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_11_port, QN => n4458);
   t_STATE_RAM0_reg_1_11_inst : FD1 port map( D => n3996, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_11_port, QN => n_3342);
   t_STATE_RAM0_reg_2_11_inst : FD1 port map( D => n3995, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_11_port, QN => n_3343);
   t_STATE_RAM0_reg_3_11_inst : FD1 port map( D => n3994, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_11_port, QN => n_3344);
   v_RAM_OUT0_reg_11_inst : FD1 port map( D => n3993, CP => CLK_I, Q => 
                           v_RAM_OUT0_11_port, QN => n4408);
   v_RAM_IN0_reg_3_inst : FD1 port map( D => n3992, CP => CLK_I, Q => 
                           v_RAM_IN0_3_port, QN => n_3345);
   t_STATE_RAM0_reg_0_3_inst : FD1 port map( D => n3991, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_3_port, QN => n4459);
   t_STATE_RAM0_reg_1_3_inst : FD1 port map( D => n3990, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_3_port, QN => n_3346);
   t_STATE_RAM0_reg_2_3_inst : FD1 port map( D => n3989, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_3_port, QN => n_3347);
   t_STATE_RAM0_reg_3_3_inst : FD1 port map( D => n3988, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_3_port, QN => n_3348);
   v_RAM_OUT0_reg_3_inst : FD1 port map( D => n3987, CP => CLK_I, Q => 
                           v_RAM_OUT0_3_port, QN => n4365);
   v_RAM_IN0_reg_8_inst : FD1 port map( D => n3986, CP => CLK_I, Q => 
                           v_RAM_IN0_8_port, QN => n_3349);
   t_STATE_RAM0_reg_0_8_inst : FD1 port map( D => n3985, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_8_port, QN => n4460);
   t_STATE_RAM0_reg_1_8_inst : FD1 port map( D => n3984, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_8_port, QN => n_3350);
   t_STATE_RAM0_reg_2_8_inst : FD1 port map( D => n3983, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_8_port, QN => n_3351);
   t_STATE_RAM0_reg_3_8_inst : FD1 port map( D => n3982, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_8_port, QN => n_3352);
   v_RAM_OUT0_reg_8_inst : FD1 port map( D => n3981, CP => CLK_I, Q => 
                           v_RAM_OUT0_8_port, QN => n4352);
   v_RAM_IN0_reg_16_inst : FD1 port map( D => n3980, CP => CLK_I, Q => 
                           v_RAM_IN0_16_port, QN => n4377);
   t_STATE_RAM0_reg_0_16_inst : FD1 port map( D => n3979, CP => CLK_I, Q => 
                           n_3353, QN => n4426);
   t_STATE_RAM0_reg_1_16_inst : FD1 port map( D => n3978, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_16_port, QN => n_3354);
   t_STATE_RAM0_reg_2_16_inst : FD1 port map( D => n3977, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_16_port, QN => n_3355);
   t_STATE_RAM0_reg_3_16_inst : FD1 port map( D => n3976, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_16_port, QN => n_3356);
   v_RAM_OUT0_reg_16_inst : FD1 port map( D => n3975, CP => CLK_I, Q => 
                           v_RAM_OUT0_16_port, QN => n4354);
   v_RAM_IN0_reg_0_inst : FD1 port map( D => n3974, CP => CLK_I, Q => 
                           v_RAM_IN0_0_port, QN => n_3357);
   t_STATE_RAM0_reg_0_0_inst : FD1 port map( D => n3973, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_0_port, QN => n4461);
   t_STATE_RAM0_reg_1_0_inst : FD1 port map( D => n3972, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_0_port, QN => n_3358);
   t_STATE_RAM0_reg_2_0_inst : FD1 port map( D => n3971, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_0_port, QN => n_3359);
   t_STATE_RAM0_reg_3_0_inst : FD1 port map( D => n3970, CP => CLK_I, Q => 
                           t_STATE_RAM0_3_0_port, QN => n_3360);
   v_RAM_OUT0_reg_0_inst : FD1 port map( D => n3969, CP => CLK_I, Q => 
                           v_RAM_OUT0_0_port, QN => n4356);
   DATA_O_reg_7_inst : FD1 port map( D => n3968, CP => CLK_I, Q => 
                           DATA_O_7_port, QN => n_3361);
   DATA_O_reg_6_inst : FD1 port map( D => n3967, CP => CLK_I, Q => 
                           DATA_O_6_port, QN => n_3362);
   DATA_O_reg_5_inst : FD1 port map( D => n3966, CP => CLK_I, Q => 
                           DATA_O_5_port, QN => n_3363);
   DATA_O_reg_4_inst : FD1 port map( D => n3965, CP => CLK_I, Q => 
                           DATA_O_4_port, QN => n_3364);
   DATA_O_reg_3_inst : FD1 port map( D => n3964, CP => CLK_I, Q => 
                           DATA_O_3_port, QN => n_3365);
   DATA_O_reg_2_inst : FD1 port map( D => n3963, CP => CLK_I, Q => 
                           DATA_O_2_port, QN => n_3366);
   DATA_O_reg_1_inst : FD1 port map( D => n3962, CP => CLK_I, Q => 
                           DATA_O_1_port, QN => n_3367);
   DATA_O_reg_0_inst : FD1 port map( D => n3961, CP => CLK_I, Q => 
                           DATA_O_0_port, QN => n_3368);
   VALID_O_reg : FD1 port map( D => n3960, CP => CLK_I, Q => VALID_O, QN => 
                           n3813);
   KEXP0 : key_expansion port map( KEY_I(7) => KEY_I(7), KEY_I(6) => KEY_I(6), 
                           KEY_I(5) => KEY_I(5), KEY_I(4) => KEY_I(4), KEY_I(3)
                           => KEY_I(3), KEY_I(2) => KEY_I(2), KEY_I(1) => 
                           KEY_I(1), KEY_I(0) => KEY_I(0), VALID_KEY_I => 
                           VALID_KEY_I, CLK_I => CLK_I, RESET_I => RESET_I, 
                           CE_I => CE_I, DONE_O => KEY_READY_O, GET_KEY_I => 
                           GET_KEY, KEY_NUMB_I(5) => v_INV_KEY_NUMB_5_port, 
                           KEY_NUMB_I(4) => v_INV_KEY_NUMB_4_port, 
                           KEY_NUMB_I(3) => v_INV_KEY_NUMB_3_port, 
                           KEY_NUMB_I(2) => v_INV_KEY_NUMB_2_port, 
                           KEY_NUMB_I(1) => n4435, KEY_NUMB_I(0) => n4419, 
                           KEY_EXP_O(31) => v_KEY_COLUMN_31_port, KEY_EXP_O(30)
                           => v_KEY_COLUMN_30_port, KEY_EXP_O(29) => 
                           v_KEY_COLUMN_29_port, KEY_EXP_O(28) => 
                           v_KEY_COLUMN_28_port, KEY_EXP_O(27) => 
                           v_KEY_COLUMN_27_port, KEY_EXP_O(26) => 
                           v_KEY_COLUMN_26_port, KEY_EXP_O(25) => 
                           v_KEY_COLUMN_25_port, KEY_EXP_O(24) => 
                           v_KEY_COLUMN_24_port, KEY_EXP_O(23) => 
                           v_KEY_COLUMN_23_port, KEY_EXP_O(22) => 
                           v_KEY_COLUMN_22_port, KEY_EXP_O(21) => 
                           v_KEY_COLUMN_21_port, KEY_EXP_O(20) => 
                           v_KEY_COLUMN_20_port, KEY_EXP_O(19) => 
                           v_KEY_COLUMN_19_port, KEY_EXP_O(18) => 
                           v_KEY_COLUMN_18_port, KEY_EXP_O(17) => 
                           v_KEY_COLUMN_17_port, KEY_EXP_O(16) => 
                           v_KEY_COLUMN_16_port, KEY_EXP_O(15) => 
                           v_KEY_COLUMN_15_port, KEY_EXP_O(14) => 
                           v_KEY_COLUMN_14_port, KEY_EXP_O(13) => 
                           v_KEY_COLUMN_13_port, KEY_EXP_O(12) => 
                           v_KEY_COLUMN_12_port, KEY_EXP_O(11) => 
                           v_KEY_COLUMN_11_port, KEY_EXP_O(10) => 
                           v_KEY_COLUMN_10_port, KEY_EXP_O(9) => 
                           v_KEY_COLUMN_9_port, KEY_EXP_O(8) => 
                           v_KEY_COLUMN_8_port, KEY_EXP_O(7) => 
                           v_KEY_COLUMN_7_port, KEY_EXP_O(6) => 
                           v_KEY_COLUMN_6_port, KEY_EXP_O(5) => 
                           v_KEY_COLUMN_5_port, KEY_EXP_O(4) => 
                           v_KEY_COLUMN_4_port, KEY_EXP_O(3) => 
                           v_KEY_COLUMN_3_port, KEY_EXP_O(2) => 
                           v_KEY_COLUMN_2_port, KEY_EXP_O(1) => 
                           v_KEY_COLUMN_1_port, KEY_EXP_O(0) => 
                           v_KEY_COLUMN_0_port);
   U4208 : MUX21H port map( A => v_DATA_COLUMN_7_port, B => DATA_I(7), S => 
                           n4492, Z => n7946);
   U4209 : MUX21H port map( A => v_DATA_COLUMN_31_port, B => DATA_I(7), S => 
                           n4493, Z => n7947);
   U4210 : MUX21H port map( A => DATA_I(7), B => v_DATA_COLUMN_23_port, S => 
                           n4494, Z => n7948);
   U4211 : MUX21H port map( A => v_DATA_COLUMN_15_port, B => DATA_I(7), S => 
                           n4495, Z => n7949);
   U4212 : MUX21H port map( A => v_DATA_COLUMN_6_port, B => DATA_I(6), S => 
                           n4492, Z => n7950);
   U4213 : MUX21H port map( A => v_DATA_COLUMN_30_port, B => DATA_I(6), S => 
                           n4493, Z => n7951);
   U4214 : MUX21H port map( A => DATA_I(6), B => v_DATA_COLUMN_22_port, S => 
                           n4494, Z => n7952);
   U4215 : MUX21H port map( A => v_DATA_COLUMN_14_port, B => DATA_I(6), S => 
                           n4495, Z => n7953);
   U4216 : MUX21H port map( A => v_DATA_COLUMN_5_port, B => DATA_I(5), S => 
                           n4492, Z => n7954);
   U4217 : MUX21H port map( A => v_DATA_COLUMN_29_port, B => DATA_I(5), S => 
                           n4493, Z => n7955);
   U4218 : MUX21H port map( A => DATA_I(5), B => v_DATA_COLUMN_21_port, S => 
                           n4494, Z => n7956);
   U4219 : MUX21H port map( A => v_DATA_COLUMN_13_port, B => DATA_I(5), S => 
                           n4495, Z => n7957);
   U4220 : MUX21H port map( A => v_DATA_COLUMN_4_port, B => DATA_I(4), S => 
                           n4492, Z => n7958);
   U4221 : MUX21H port map( A => v_DATA_COLUMN_28_port, B => DATA_I(4), S => 
                           n4493, Z => n7959);
   U4222 : MUX21H port map( A => DATA_I(4), B => v_DATA_COLUMN_20_port, S => 
                           n4494, Z => n7960);
   U4223 : MUX21H port map( A => v_DATA_COLUMN_12_port, B => DATA_I(4), S => 
                           n4495, Z => n7961);
   U4224 : MUX21H port map( A => v_DATA_COLUMN_3_port, B => DATA_I(3), S => 
                           n4492, Z => n7962);
   U4225 : MUX21H port map( A => v_DATA_COLUMN_27_port, B => DATA_I(3), S => 
                           n4493, Z => n7963);
   U4226 : MUX21H port map( A => DATA_I(3), B => v_DATA_COLUMN_19_port, S => 
                           n4494, Z => n7964);
   U4227 : MUX21H port map( A => v_DATA_COLUMN_11_port, B => DATA_I(3), S => 
                           n4495, Z => n7965);
   U4228 : MUX21H port map( A => v_DATA_COLUMN_2_port, B => DATA_I(2), S => 
                           n4492, Z => n7966);
   U4229 : MUX21H port map( A => v_DATA_COLUMN_26_port, B => DATA_I(2), S => 
                           n4493, Z => n7967);
   U4230 : MUX21H port map( A => DATA_I(2), B => v_DATA_COLUMN_18_port, S => 
                           n4494, Z => n7968);
   U4231 : MUX21H port map( A => v_DATA_COLUMN_10_port, B => DATA_I(2), S => 
                           n4495, Z => n7969);
   U4232 : MUX21H port map( A => v_DATA_COLUMN_9_port, B => DATA_I(1), S => 
                           n4495, Z => n7970);
   U4233 : MUX21H port map( A => v_DATA_COLUMN_25_port, B => DATA_I(1), S => 
                           n4493, Z => n7971);
   U4234 : MUX21H port map( A => v_DATA_COLUMN_1_port, B => DATA_I(1), S => 
                           n4492, Z => n7972);
   U4235 : MUX21H port map( A => DATA_I(1), B => v_DATA_COLUMN_17_port, S => 
                           n4494, Z => n7973);
   U4236 : AO1 port map( A => n4414, B => n4496, C => n4497, D => n4498, Z => 
                           n7974);
   U4237 : MUX21L port map( A => n4499, B => n4500, S => 
                           v_CALCULATION_CNTR_7_port, Z => n7975);
   U4238 : AO6 port map( A => n4501, B => n4417, C => n4502, Z => n4500);
   U4239 : ND2 port map( A => v_CALCULATION_CNTR_6_port, B => n4503, Z => n4499
                           );
   U4240 : MUX21H port map( A => n4502, B => n4503, S => n4417, Z => n7976);
   U4241 : AN3 port map( A => n4501, B => n4504, C => v_CALCULATION_CNTR_5_port
                           , Z => n4503);
   U4242 : AO7 port map( A => v_CALCULATION_CNTR_5_port, B => n4505, C => n4506
                           , Z => n4502);
   U4243 : MUX21L port map( A => n4507, B => n4506, S => 
                           v_CALCULATION_CNTR_5_port, Z => n7977);
   U4244 : AO6 port map( A => n4508, B => n4501, C => n4509, Z => n4506);
   U4245 : IV port map( A => n4504, Z => n4508);
   U4246 : ND2 port map( A => n4501, B => n4504, Z => n4507);
   U4247 : AN3 port map( A => v_CALCULATION_CNTR_3_port, B => 
                           v_CALCULATION_CNTR_4_port, C => n4510, Z => n4504);
   U4248 : MUX21L port map( A => CE_I, B => n4511, S => n4418, Z => n4349);
   U4249 : MUX21H port map( A => v_DATA_COLUMN_24_port, B => DATA_I(0), S => 
                           n4493, Z => n4348);
   U4250 : AN3 port map( A => v_CNT4_0_port, B => VALID_DATA_I, C => 
                           v_CNT4_1_port, Z => n4493);
   U4251 : ND2 port map( A => n4512, B => n4494, Z => n4340);
   U4252 : MUX21L port map( A => n4495, B => v_CNT4_1_port, S => n4513, Z => 
                           n4512);
   U4253 : MUX21H port map( A => v_DATA_COLUMN_8_port, B => DATA_I(0), S => 
                           n4495, Z => n4339);
   U4254 : AN3 port map( A => VALID_DATA_I, B => n4370, C => v_CNT4_0_port, Z 
                           => n4495);
   U4255 : MUX21H port map( A => DATA_I(0), B => v_DATA_COLUMN_16_port, S => 
                           n4494, Z => n4331);
   U4256 : MUX21H port map( A => v_DATA_COLUMN_0_port, B => DATA_I(0), S => 
                           n4492, Z => n4323);
   U4257 : AN3 port map( A => n4418, B => n4370, C => VALID_DATA_I, Z => n4492)
                           ;
   U4258 : AO4 port map( A => RESET_I, B => n4511, C => n4514, D => n4432, Z =>
                           n4315);
   U4259 : NR2 port map( A => RESET_I, B => n4513, Z => n4514);
   U4260 : AO4 port map( A => n4515, B => n4400, C => n4516, D => n4517, Z => 
                           n4314);
   U4261 : ND3 port map( A => n4518, B => n7894, C => n7893, Z => n4517);
   U4262 : ND4 port map( A => n4519, B => CE_I, C => v_CALCULATION_CNTR_0_port,
                           D => n4369, Z => n4516);
   U4263 : NR2 port map( A => n4509, B => n4520, Z => n4515);
   U4264 : MUX21L port map( A => n4521, B => n4505, S => n4399, Z => n4313);
   U4265 : MUX21L port map( A => n4522, B => n4523, S => n4405, Z => n4312);
   U4266 : ND2 port map( A => n4501, B => v_CALCULATION_CNTR_0_port, Z => n4523
                           );
   U4267 : AO6 port map( A => n4501, B => n4399, C => n4509, Z => n4522);
   U4268 : IV port map( A => n4524, Z => n4311);
   U4269 : AO2 port map( A => v_CALCULATION_CNTR_2_port, B => n4509, C => n4525
                           , D => n4501, Z => n4524);
   U4270 : ND2 port map( A => n4526, B => n4527, Z => n4525);
   U4271 : MUX21L port map( A => n4528, B => v_CALCULATION_CNTR_2_port, S => 
                           n4405, Z => n4527);
   U4272 : MUX21L port map( A => n4529, B => n4530, S => n4401, Z => n4310);
   U4273 : ND2 port map( A => n4501, B => n4510, Z => n4530);
   U4274 : IV port map( A => n4505, Z => n4501);
   U4275 : AO4 port map( A => n4529, B => n4416, C => n4531, D => n4505, Z => 
                           n4309);
   U4276 : AO6 port map( A => n4532, B => n4510, C => n4533, Z => n4531);
   U4277 : NR2 port map( A => v_CALCULATION_CNTR_4_port, B => n4401, Z => n4532
                           );
   U4278 : IV port map( A => n4534, Z => n4529);
   U4279 : AO7 port map( A => n4510, B => n4505, C => n4521, Z => n4534);
   U4280 : ND3 port map( A => n4535, B => n4521, C => n4520, Z => n4505);
   U4281 : NR2 port map( A => n4536, B => n4405, Z => n4510);
   U4282 : MUX21H port map( A => n7896, B => GET_KEY, S => CE_I, Z => n4305);
   U4283 : MUX21H port map( A => n7891, B => n7896, S => CE_I, Z => n4304);
   U4284 : AO1 port map( A => n4433, B => n4537, C => n4497, D => n4538, Z => 
                           n4303);
   U4285 : IV port map( A => n4496, Z => n4538);
   U4286 : ND2 port map( A => n7891, B => CE_I, Z => n4537);
   U4287 : ND2 port map( A => n4539, B => n4540, Z => n4301);
   U4288 : EO port map( A => n4541, B => n3947, Z => n4539);
   U4289 : NR2 port map( A => v_INV_KEY_NUMB_4_port, B => n4542, Z => n4541);
   U4290 : ND2 port map( A => n4543, B => n4540, Z => n4300);
   U4291 : EN port map( A => n4419, B => n4544, Z => n4543);
   U4292 : AO3 port map( A => n4544, B => n4545, C => n4546, D => n4540, Z => 
                           n4299);
   U4293 : AO7 port map( A => n4544, B => v_KEY_NUMB_0_port, C => 
                           v_KEY_NUMB_1_port, Z => n4546);
   U4294 : IV port map( A => n4547, Z => n4545);
   U4295 : MUX21L port map( A => n4411, B => n4548, S => n4549, Z => n4298);
   U4296 : AO3 port map( A => n7886, B => n4550, C => n4551, D => n4552, Z => 
                           n4548);
   U4297 : AO7 port map( A => n4547, B => n4411, C => n4553, Z => n4551);
   U4298 : AO3 port map( A => n4554, B => n4429, C => n4542, D => n4540, Z => 
                           n4297);
   U4299 : ND2 port map( A => n4555, B => n4540, Z => n4296);
   U4300 : ND2 port map( A => n4549, B => n4556, Z => n4540);
   U4301 : AO7 port map( A => n7886, B => n4550, C => n4552, Z => n4556);
   U4302 : IV port map( A => n4544, Z => n4549);
   U4303 : EO port map( A => v_INV_KEY_NUMB_4_port, B => n4542, Z => n4555);
   U4304 : ND2 port map( A => n4554, B => n4429, Z => n4542);
   U4305 : NR2 port map( A => n4553, B => n4544, Z => n4554);
   U4306 : AO6 port map( A => GET_KEY, B => CE_I, C => n4497, Z => n4544);
   U4307 : AO7 port map( A => n7886, B => n4511, C => n4552, Z => n4497);
   U4308 : ND2 port map( A => CE_I, B => VALID_DATA_I, Z => n4511);
   U4309 : ND2 port map( A => n4547, B => n4411, Z => n4553);
   U4310 : NR2 port map( A => v_KEY_NUMB_0_port, B => v_KEY_NUMB_1_port, Z => 
                           n4547);
   U4311 : AO4 port map( A => n4557, B => n4434, C => n4558, D => n4559, Z => 
                           n4295);
   U4312 : ND2 port map( A => n4560, B => n4561, Z => n4559);
   U4313 : AO7 port map( A => n4557, B => n4415, C => n4562, Z => n4294);
   U4314 : AO3 port map( A => n4563, B => n4564, C => n4561, D => n4560, Z => 
                           n4562);
   U4315 : AO7 port map( A => n4399, B => n4565, C => n4566, Z => n4561);
   U4316 : NR2 port map( A => n4509, B => n4567, Z => n4557);
   U4317 : AO6 port map( A => n4568, B => n4560, C => RESET_I, Z => n4567);
   U4318 : IV port map( A => n4565, Z => n4568);
   U4319 : AO3 port map( A => n4431, B => n4521, C => n4569, D => n4570, Z => 
                           n4293);
   U4320 : ND4 port map( A => n7886, B => CE_I, C => n4552, D => n4550, Z => 
                           n4570);
   U4321 : AO7 port map( A => n4571, B => n4400, C => n4520, Z => n4569);
   U4322 : IV port map( A => n4509, Z => n4521);
   U4323 : NR2 port map( A => RESET_I, B => CE_I, Z => n4509);
   U4324 : MUX21H port map( A => n4518, B => n7895, S => n4572, Z => n4292);
   U4325 : MUX21L port map( A => n4573, B => n4574, S => n7892, Z => n4291);
   U4326 : MUX21H port map( A => n4575, B => n4576, S => n7893, Z => n4290);
   U4327 : NR2 port map( A => n4573, B => n4369, Z => n4575);
   U4328 : MUX21L port map( A => n4577, B => n4578, S => n7894, Z => n4289);
   U4329 : AO6 port map( A => n4520, B => n4430, C => n4576, Z => n4578);
   U4330 : AO7 port map( A => n7892, B => n4579, C => n4574, Z => n4576);
   U4331 : NR2 port map( A => n4572, B => n4518, Z => n4574);
   U4332 : NR2 port map( A => n4579, B => n7895, Z => n4518);
   U4333 : OR3 port map( A => n4369, B => n4430, C => n4573, Z => n4577);
   U4334 : OR3 port map( A => n4579, B => n4572, C => n4436, Z => n4573);
   U4335 : NR2 port map( A => RESET_I, B => n4580, Z => n4572);
   U4336 : AO6 port map( A => n7945, B => n4535, C => n4513, Z => n4580);
   U4337 : MUX21L port map( A => n4581, B => n4582, S => n4400, Z => n4535);
   U4338 : AN2 port map( A => v_CALCULATION_CNTR_0_port, B => n4519, Z => n4582
                           );
   U4339 : IV port map( A => n4520, Z => n4579);
   U4340 : NR2 port map( A => n4431, B => RESET_I, Z => n4520);
   U4341 : AO7 port map( A => n4583, B => n4584, C => n4585, Z => n4288);
   U4342 : AO2 port map( A => n4586, B => n4587, C => n7851, D => n4588, Z => 
                           n4585);
   U4343 : AO7 port map( A => n4589, B => n4584, C => n4590, Z => n4287);
   U4344 : AO2 port map( A => n4591, B => n4587, C => n7850, D => n4588, Z => 
                           n4590);
   U4345 : AO7 port map( A => n4592, B => n4584, C => n4593, Z => n4286);
   U4346 : AO2 port map( A => n4587, B => n4594, C => n7849, D => n4588, Z => 
                           n4593);
   U4347 : AO7 port map( A => n4595, B => n4584, C => n4596, Z => n4285);
   U4348 : AO2 port map( A => n4597, B => n4587, C => n7852, D => n4588, Z => 
                           n4596);
   U4349 : AO7 port map( A => n4598, B => n4584, C => n4599, Z => n4284);
   U4350 : AO2 port map( A => n4600, B => n4587, C => n7859, D => n4588, Z => 
                           n4599);
   U4351 : AO7 port map( A => n4601, B => n4584, C => n4602, Z => n4283);
   U4352 : AO2 port map( A => n4603, B => n4587, C => n7867, D => n4588, Z => 
                           n4602);
   U4353 : AO7 port map( A => n4604, B => n4584, C => n4605, Z => n4282);
   U4354 : AO2 port map( A => n4606, B => n4587, C => n7853, D => n4588, Z => 
                           n4605);
   U4355 : AO7 port map( A => n4607, B => n4584, C => n4608, Z => n4281);
   U4356 : AO2 port map( A => n4609, B => n4587, C => n7858, D => n4588, Z => 
                           n4608);
   U4357 : NR2 port map( A => n4610, B => n4588, Z => n4587);
   U4358 : NR2 port map( A => n4610, B => n4611, Z => n4588);
   U4359 : IV port map( A => n4612, Z => n4607);
   U4360 : AO7 port map( A => n4613, B => n4584, C => n4614, Z => n4280);
   U4361 : AO2 port map( A => n4615, B => n4616, C => n7848, D => n4617, Z => 
                           n4614);
   U4362 : AO7 port map( A => n4618, B => n4584, C => n4619, Z => n4279);
   U4363 : AO2 port map( A => n4620, B => n4616, C => n7847, D => n4617, Z => 
                           n4619);
   U4364 : IV port map( A => n4621, Z => n4618);
   U4365 : AO7 port map( A => n4622, B => n4584, C => n4623, Z => n4278);
   U4366 : AO2 port map( A => n4624, B => n4616, C => n7877, D => n4617, Z => 
                           n4623);
   U4367 : AO7 port map( A => n4625, B => n4584, C => n4626, Z => n4277);
   U4368 : AO2 port map( A => n4627, B => n4616, C => n7846, D => n4617, Z => 
                           n4626);
   U4369 : AO7 port map( A => n4628, B => n4584, C => n4629, Z => n4276);
   U4370 : AO2 port map( A => n4630, B => n4616, C => n7845, D => n4617, Z => 
                           n4629);
   U4371 : AO7 port map( A => n4631, B => n4584, C => n4632, Z => n4275);
   U4372 : AO2 port map( A => n4616, B => n4633, C => n7844, D => n4617, Z => 
                           n4632);
   U4373 : AO7 port map( A => n4361, B => n4634, C => n4635, Z => n4633);
   U4374 : AO2 port map( A => n4636, B => n4637, C => n4638, D => n4639, Z => 
                           n4635);
   U4375 : AO1 port map( A => v_RAM_OUT0_13_port, B => n4640, C => n4641, D => 
                           n4642, Z => n4637);
   U4376 : NR2 port map( A => n4643, B => n4644, Z => n4641);
   U4377 : AO1 port map( A => n4645, B => n4646, C => n4647, D => n4648, Z => 
                           n4636);
   U4378 : NR2 port map( A => n4649, B => n4650, Z => n4648);
   U4379 : IV port map( A => n4651, Z => n4650);
   U4380 : AO7 port map( A => n4652, B => n4584, C => n4653, Z => n4274);
   U4381 : AO2 port map( A => n4654, B => n4616, C => n7866, D => n4617, Z => 
                           n4653);
   U4382 : AO7 port map( A => n4655, B => n4584, C => n4656, Z => n4273);
   U4383 : AO2 port map( A => n4657, B => n4616, C => n7876, D => n4617, Z => 
                           n4656);
   U4384 : NR2 port map( A => n4610, B => n4617, Z => n4616);
   U4385 : NR2 port map( A => n4610, B => n4658, Z => n4617);
   U4386 : MUX21L port map( A => n4659, B => n4660, S => n4361, Z => n4657);
   U4387 : AO3 port map( A => n4661, B => n4662, C => n4663, D => n4664, Z => 
                           n4659);
   U4388 : AO2 port map( A => n4665, B => n4666, C => n4667, D => n4668, Z => 
                           n4664);
   U4389 : ND3 port map( A => v_RAM_OUT0_15_port, B => n4353, C => n4669, Z => 
                           n4663);
   U4390 : MUX21L port map( A => n4670, B => n4671, S => n4672, Z => n4669);
   U4391 : MUX21L port map( A => n4673, B => n4674, S => n4357, Z => n4670);
   U4392 : MUX21L port map( A => n4675, B => n4676, S => n4672, Z => n4662);
   U4393 : MUX21L port map( A => n4677, B => n4678, S => n4357, Z => n4675);
   U4394 : AO7 port map( A => n4679, B => n4584, C => n4680, Z => n4272);
   U4395 : AO2 port map( A => n4681, B => n4682, C => n7897, D => n4683, Z => 
                           n4680);
   U4396 : AO7 port map( A => n4684, B => n4584, C => n4685, Z => n4271);
   U4397 : AO2 port map( A => n4686, B => n4682, C => n7903, D => n4683, Z => 
                           n4685);
   U4398 : AO7 port map( A => n4687, B => n4584, C => n4688, Z => n4270);
   U4399 : AO2 port map( A => n4682, B => n4689, C => n7909, D => n4683, Z => 
                           n4688);
   U4400 : IV port map( A => n4690, Z => n4687);
   U4401 : AO7 port map( A => n4691, B => n4584, C => n4692, Z => n4269);
   U4402 : AO2 port map( A => n4693, B => n4682, C => n7915, D => n4683, Z => 
                           n4692);
   U4403 : AO7 port map( A => n4694, B => n4584, C => n4695, Z => n4268);
   U4404 : AO2 port map( A => n4696, B => n4682, C => n7921, D => n4683, Z => 
                           n4695);
   U4405 : AO7 port map( A => n4697, B => n4584, C => n4698, Z => n4267);
   U4406 : AO2 port map( A => n4699, B => n4682, C => n7927, D => n4683, Z => 
                           n4698);
   U4407 : AO7 port map( A => n4700, B => n4584, C => n4701, Z => n4266);
   U4408 : AO2 port map( A => n4702, B => n4682, C => n7933, D => n4683, Z => 
                           n4701);
   U4409 : AO7 port map( A => n4703, B => n4584, C => n4704, Z => n4265);
   U4410 : AO2 port map( A => n4705, B => n4682, C => n7939, D => n4683, Z => 
                           n4704);
   U4411 : NR2 port map( A => n4610, B => n4683, Z => n4682);
   U4412 : NR2 port map( A => n4610, B => n4706, Z => n4683);
   U4413 : AO7 port map( A => n4707, B => n4584, C => n4708, Z => n4264);
   U4414 : AO2 port map( A => n4709, B => n4710, C => n7898, D => n4711, Z => 
                           n4708);
   U4415 : AO7 port map( A => n4712, B => n4584, C => n4713, Z => n4263);
   U4416 : AO2 port map( A => n4714, B => n4710, C => n7904, D => n4711, Z => 
                           n4713);
   U4417 : AO7 port map( A => n4715, B => n4584, C => n4716, Z => n4262);
   U4418 : AO2 port map( A => n4710, B => n4717, C => n7910, D => n4711, Z => 
                           n4716);
   U4419 : AO7 port map( A => n4718, B => n4584, C => n4719, Z => n4261);
   U4420 : AO2 port map( A => n4720, B => n4710, C => n7916, D => n4711, Z => 
                           n4719);
   U4421 : AO7 port map( A => n4721, B => n4584, C => n4722, Z => n4260);
   U4422 : AO2 port map( A => n4723, B => n4710, C => n7922, D => n4711, Z => 
                           n4722);
   U4423 : AO7 port map( A => n4724, B => n4584, C => n4725, Z => n4259);
   U4424 : AO2 port map( A => n4726, B => n4710, C => n7928, D => n4711, Z => 
                           n4725);
   U4425 : AO7 port map( A => n4727, B => n4584, C => n4728, Z => n4258);
   U4426 : AO2 port map( A => n4729, B => n4710, C => n7934, D => n4711, Z => 
                           n4728);
   U4427 : AO7 port map( A => n4730, B => n4584, C => n4731, Z => n4257);
   U4428 : AO2 port map( A => n4732, B => n4710, C => n7940, D => n4711, Z => 
                           n4731);
   U4429 : NR2 port map( A => n4610, B => n4711, Z => n4710);
   U4430 : NR2 port map( A => n4610, B => n4733, Z => n4711);
   U4431 : AO7 port map( A => n4734, B => n4735, C => n4736, Z => n4256);
   U4432 : AO2 port map( A => n4737, B => n4586, C => n7899, D => n4738, Z => 
                           n4736);
   U4433 : AO7 port map( A => n4739, B => n4735, C => n4740, Z => n4255);
   U4434 : AO2 port map( A => n4737, B => n4591, C => n7905, D => n4738, Z => 
                           n4740);
   U4435 : AO7 port map( A => n4741, B => n4735, C => n4742, Z => n4254);
   U4436 : AO2 port map( A => n4737, B => n4594, C => n7911, D => n4738, Z => 
                           n4742);
   U4437 : AO7 port map( A => n4743, B => n4735, C => n4744, Z => n4253);
   U4438 : AO2 port map( A => n4737, B => n4597, C => n7917, D => n4738, Z => 
                           n4744);
   U4439 : AO7 port map( A => n4745, B => n4735, C => n4746, Z => n4252);
   U4440 : AO2 port map( A => n4737, B => n4600, C => n7923, D => n4738, Z => 
                           n4746);
   U4441 : AO7 port map( A => n4747, B => n4735, C => n4748, Z => n4251);
   U4442 : AO2 port map( A => n4737, B => n4603, C => n7929, D => n4738, Z => 
                           n4748);
   U4443 : AO7 port map( A => n4749, B => n4735, C => n4750, Z => n4250);
   U4444 : AO2 port map( A => n4737, B => n4606, C => n7935, D => n4738, Z => 
                           n4750);
   U4445 : AO7 port map( A => n4751, B => n4735, C => n4752, Z => n4249);
   U4446 : AO2 port map( A => n4737, B => n4609, C => n7941, D => n4738, Z => 
                           n4752);
   U4447 : NR2 port map( A => n4753, B => n4738, Z => n4737);
   U4448 : NR2 port map( A => n4753, B => n4733, Z => n4738);
   U4449 : AO7 port map( A => n4754, B => n4735, C => n4755, Z => n4248);
   U4450 : AO2 port map( A => n4756, B => n4615, C => n7843, D => n4757, Z => 
                           n4755);
   U4451 : AO7 port map( A => n4758, B => n4735, C => n4759, Z => n4247);
   U4452 : AO2 port map( A => n4756, B => n4620, C => n7842, D => n4757, Z => 
                           n4759);
   U4453 : IV port map( A => n4760, Z => n4758);
   U4454 : AO7 port map( A => n4761, B => n4735, C => n4762, Z => n4246);
   U4455 : AO2 port map( A => n4756, B => n4624, C => n7880, D => n4757, Z => 
                           n4762);
   U4456 : AO7 port map( A => n4763, B => n4735, C => n4764, Z => n4245);
   U4457 : AO2 port map( A => n4756, B => n4627, C => n7841, D => n4757, Z => 
                           n4764);
   U4458 : AO7 port map( A => n4765, B => n4735, C => n4766, Z => n4244);
   U4459 : AO2 port map( A => n4756, B => n4630, C => n7840, D => n4757, Z => 
                           n4766);
   U4460 : AO7 port map( A => n4767, B => n4735, C => n4768, Z => n4243);
   U4461 : AO2 port map( A => n4769, B => n4756, C => n7839, D => n4757, Z => 
                           n4768);
   U4462 : AO7 port map( A => n4770, B => n4735, C => n4771, Z => n4242);
   U4463 : AO2 port map( A => n4756, B => n4654, C => n7838, D => n4757, Z => 
                           n4771);
   U4464 : AO7 port map( A => n4772, B => n4735, C => n4773, Z => n4241);
   U4465 : AO2 port map( A => n4774, B => n4756, C => n7879, D => n4757, Z => 
                           n4773);
   U4466 : NR2 port map( A => n4753, B => n4757, Z => n4756);
   U4467 : NR2 port map( A => n4753, B => n4611, Z => n4757);
   U4468 : AO7 port map( A => n4775, B => n4735, C => n4776, Z => n4240);
   U4469 : AO2 port map( A => n4777, B => n4681, C => n7837, D => n4778, Z => 
                           n4776);
   U4470 : AO7 port map( A => n4779, B => n4735, C => n4780, Z => n4239);
   U4471 : AO2 port map( A => n4777, B => n4686, C => n7836, D => n4778, Z => 
                           n4780);
   U4472 : AO7 port map( A => n4781, B => n4735, C => n4782, Z => n4238);
   U4473 : AO2 port map( A => n4777, B => n4689, C => n7835, D => n4778, Z => 
                           n4782);
   U4474 : IV port map( A => n4783, Z => n4781);
   U4475 : AO7 port map( A => n4784, B => n4735, C => n4785, Z => n4237);
   U4476 : AO2 port map( A => n4777, B => n4693, C => n7834, D => n4778, Z => 
                           n4785);
   U4477 : AO7 port map( A => n4786, B => n4735, C => n4787, Z => n4236);
   U4478 : AO2 port map( A => n4777, B => n4696, C => n7864, D => n4778, Z => 
                           n4787);
   U4479 : AO7 port map( A => n4788, B => n4735, C => n4789, Z => n4235);
   U4480 : AO2 port map( A => n4790, B => n4777, C => n7872, D => n4778, Z => 
                           n4789);
   U4481 : MUX21L port map( A => n4791, B => n4792, S => n4395, Z => n4790);
   U4482 : AO1 port map( A => n4793, B => n4794, C => n4795, D => n4796, Z => 
                           n4791);
   U4483 : AO4 port map( A => n4797, B => n4798, C => n4799, D => n4800, Z => 
                           n4796);
   U4484 : AO6 port map( A => n4801, B => n4802, C => n4803, Z => n4799);
   U4485 : AO4 port map( A => n4358, B => n4804, C => n4805, D => n4806, Z => 
                           n4803);
   U4486 : AO4 port map( A => n4403, B => n4807, C => n4808, D => n4809, Z => 
                           n4795);
   U4487 : AO7 port map( A => n4810, B => n4735, C => n4811, Z => n4234);
   U4488 : AO2 port map( A => n4777, B => n4702, C => n7833, D => n4778, Z => 
                           n4811);
   U4489 : AO7 port map( A => n4812, B => n4735, C => n4813, Z => n4233);
   U4490 : AO2 port map( A => n4814, B => n4777, C => n7878, D => n4778, Z => 
                           n4813);
   U4491 : NR2 port map( A => n4753, B => n4778, Z => n4777);
   U4492 : NR2 port map( A => n4753, B => n4658, Z => n4778);
   U4493 : MUX21L port map( A => n4815, B => n4816, S => n4395, Z => n4814);
   U4494 : NR2 port map( A => n4817, B => n4818, Z => n4816);
   U4495 : AN3 port map( A => n4819, B => n4820, C => n4821, Z => n4817);
   U4496 : MUX21L port map( A => n4822, B => n4823, S => n4358, Z => n4821);
   U4497 : AO6 port map( A => n4824, B => v_RAM_OUT0_21_port, C => n4825, Z => 
                           n4815);
   U4498 : AO4 port map( A => n4800, B => n4826, C => n4808, D => n4827, Z => 
                           n4825);
   U4499 : MUX21L port map( A => n4828, B => n4829, S => n4830, Z => n4827);
   U4500 : MUX21L port map( A => n4831, B => n4832, S => n4358, Z => n4828);
   U4501 : IV port map( A => n4833, Z => n4824);
   U4502 : AO7 port map( A => n4834, B => n4735, C => n4835, Z => n4232);
   U4503 : AO2 port map( A => n4836, B => n4709, C => n7832, D => n4837, Z => 
                           n4835);
   U4504 : AO7 port map( A => n4838, B => n4735, C => n4839, Z => n4231);
   U4505 : AO2 port map( A => n4836, B => n4714, C => n7831, D => n4837, Z => 
                           n4839);
   U4506 : AO7 port map( A => n4840, B => n4735, C => n4841, Z => n4230);
   U4507 : AO2 port map( A => n4836, B => n4717, C => n7830, D => n4837, Z => 
                           n4841);
   U4508 : AO7 port map( A => n4842, B => n4735, C => n4843, Z => n4229);
   U4509 : AO2 port map( A => n4836, B => n4720, C => n7857, D => n4837, Z => 
                           n4843);
   U4510 : AO7 port map( A => n4844, B => n4735, C => n4845, Z => n4228);
   U4511 : AO2 port map( A => n4836, B => n4723, C => n7829, D => n4837, Z => 
                           n4845);
   U4512 : AO7 port map( A => n4846, B => n4735, C => n4847, Z => n4227);
   U4513 : AO2 port map( A => n4836, B => n4726, C => n7871, D => n4837, Z => 
                           n4847);
   U4514 : AO7 port map( A => n4848, B => n4735, C => n4849, Z => n4226);
   U4515 : AO2 port map( A => n4836, B => n4729, C => n7863, D => n4837, Z => 
                           n4849);
   U4516 : AO7 port map( A => n4850, B => n4735, C => n4851, Z => n4225);
   U4517 : AO2 port map( A => n4836, B => n4732, C => n7828, D => n4837, Z => 
                           n4851);
   U4518 : NR2 port map( A => n4753, B => n4837, Z => n4836);
   U4519 : NR2 port map( A => n4753, B => n4706, Z => n4837);
   U4520 : AO7 port map( A => n4852, B => n4853, C => n4854, Z => n4224);
   U4521 : AO2 port map( A => n4855, B => n4586, C => n7827, D => n4856, Z => 
                           n4854);
   U4522 : AO7 port map( A => n4857, B => n4853, C => n4858, Z => n4223);
   U4523 : AO2 port map( A => n4855, B => n4591, C => n7826, D => n4856, Z => 
                           n4858);
   U4524 : AO7 port map( A => n4859, B => n4853, C => n4860, Z => n4222);
   U4525 : AO2 port map( A => n4855, B => n4594, C => n7825, D => n4856, Z => 
                           n4860);
   U4526 : AO7 port map( A => n4861, B => n4853, C => n4862, Z => n4221);
   U4527 : AO2 port map( A => n4855, B => n4597, C => n7854, D => n4856, Z => 
                           n4862);
   U4528 : AO7 port map( A => n4863, B => n4853, C => n4864, Z => n4220);
   U4529 : AO2 port map( A => n4855, B => n4600, C => n7862, D => n4856, Z => 
                           n4864);
   U4530 : AO7 port map( A => n4865, B => n4853, C => n4866, Z => n4219);
   U4531 : AO2 port map( A => n4855, B => n4603, C => n7870, D => n4856, Z => 
                           n4866);
   U4532 : MUX21L port map( A => n4867, B => n4868, S => n4394, Z => n4603);
   U4533 : AO3 port map( A => n4869, B => n4870, C => n4871, D => n4872, Z => 
                           n4867);
   U4534 : AO2 port map( A => n4873, B => n4874, C => v_RAM_OUT0_5_port, D => 
                           n4875, Z => n4872);
   U4535 : AO2 port map( A => n4876, B => n4877, C => n4878, D => n4879, Z => 
                           n4871);
   U4536 : AO3 port map( A => n4880, B => n4881, C => n4882, D => n4883, Z => 
                           n4879);
   U4537 : ND2 port map( A => n4884, B => n4885, Z => n4882);
   U4538 : ND2 port map( A => n4886, B => n4887, Z => n4877);
   U4539 : AO7 port map( A => n4888, B => n4853, C => n4889, Z => n4218);
   U4540 : AO2 port map( A => n4855, B => n4606, C => n7855, D => n4856, Z => 
                           n4889);
   U4541 : AO7 port map( A => n4890, B => n4853, C => n4891, Z => n4217);
   U4542 : AO2 port map( A => n4855, B => n4609, C => n7861, D => n4856, Z => 
                           n4891);
   U4543 : MUX21L port map( A => n4892, B => n4893, S => n4394, Z => n4609);
   U4544 : AO6 port map( A => v_RAM_OUT0_5_port, B => n4894, C => n4895, Z => 
                           n4893);
   U4545 : AO4 port map( A => n4896, B => n4897, C => n4898, D => n4899, Z => 
                           n4894);
   U4546 : AO3 port map( A => n4900, B => n4901, C => n4902, D => n4903, Z => 
                           n4892);
   U4547 : AO2 port map( A => n4878, B => n4904, C => v_RAM_OUT0_5_port, D => 
                           n4905, Z => n4903);
   U4548 : AO2 port map( A => n4906, B => n4873, C => n4907, D => n4908, Z => 
                           n4902);
   U4549 : NR2 port map( A => n4909, B => n4910, Z => n4906);
   U4550 : NR2 port map( A => n4911, B => n4856, Z => n4855);
   U4551 : NR2 port map( A => n4911, B => n4706, Z => n4856);
   U4552 : AO7 port map( A => n4912, B => n4853, C => n4913, Z => n4216);
   U4553 : AO2 port map( A => n4914, B => n4615, C => n7824, D => n4915, Z => 
                           n4913);
   U4554 : AO7 port map( A => n4916, B => n4853, C => n4917, Z => n4215);
   U4555 : AO2 port map( A => n4914, B => n4620, C => n7823, D => n4915, Z => 
                           n4917);
   U4556 : IV port map( A => n4918, Z => n4916);
   U4557 : AO7 port map( A => n4919, B => n4853, C => n4920, Z => n4214);
   U4558 : AO2 port map( A => n4914, B => n4624, C => n7882, D => n4915, Z => 
                           n4920);
   U4559 : AO7 port map( A => n4921, B => n4853, C => n4922, Z => n4213);
   U4560 : AO2 port map( A => n4914, B => n4627, C => n7822, D => n4915, Z => 
                           n4922);
   U4561 : AO7 port map( A => n4923, B => n4853, C => n4924, Z => n4212);
   U4562 : AO2 port map( A => n4914, B => n4630, C => n7821, D => n4915, Z => 
                           n4924);
   U4563 : AO7 port map( A => n4925, B => n4853, C => n4926, Z => n4211);
   U4564 : AO2 port map( A => n4914, B => n4769, C => n7820, D => n4915, Z => 
                           n4926);
   U4565 : AO7 port map( A => n4927, B => n4853, C => n4928, Z => n4210);
   U4566 : AO2 port map( A => n4914, B => n4654, C => n7868, D => n4915, Z => 
                           n4928);
   U4567 : AO7 port map( A => n4929, B => n4853, C => n4930, Z => n4209);
   U4568 : AO2 port map( A => n4914, B => n4774, C => n7881, D => n4915, Z => 
                           n4930);
   U4569 : NR2 port map( A => n4911, B => n4915, Z => n4914);
   U4570 : NR2 port map( A => n4911, B => n4733, Z => n4915);
   U4571 : AO7 port map( A => n4931, B => n4853, C => n4932, Z => n4208);
   U4572 : AO2 port map( A => n4933, B => n4681, C => n7901, D => n4934, Z => 
                           n4932);
   U4573 : AO7 port map( A => n4935, B => n4853, C => n4936, Z => n4207);
   U4574 : AO2 port map( A => n4933, B => n4686, C => n7907, D => n4934, Z => 
                           n4936);
   U4575 : AO7 port map( A => n4937, B => n4853, C => n4938, Z => n4206);
   U4576 : AO2 port map( A => n4933, B => n4689, C => n7913, D => n4934, Z => 
                           n4938);
   U4577 : IV port map( A => n4939, Z => n4937);
   U4578 : AO7 port map( A => n4940, B => n4853, C => n4941, Z => n4205);
   U4579 : AO2 port map( A => n4933, B => n4693, C => n7919, D => n4934, Z => 
                           n4941);
   U4580 : AO7 port map( A => n4942, B => n4853, C => n4943, Z => n4204);
   U4581 : AO2 port map( A => n4933, B => n4696, C => n7925, D => n4934, Z => 
                           n4943);
   U4582 : AO7 port map( A => n4944, B => n4853, C => n4945, Z => n4203);
   U4583 : AO2 port map( A => n4933, B => n4699, C => n7931, D => n4934, Z => 
                           n4945);
   U4584 : AO7 port map( A => n4946, B => n4853, C => n4947, Z => n4202);
   U4585 : AO2 port map( A => n4933, B => n4702, C => n7937, D => n4934, Z => 
                           n4947);
   U4586 : AO7 port map( A => n4948, B => n4853, C => n4949, Z => n4201);
   U4587 : AO2 port map( A => n4933, B => n4705, C => n7943, D => n4934, Z => 
                           n4949);
   U4588 : NR2 port map( A => n4911, B => n4934, Z => n4933);
   U4589 : NR2 port map( A => n4911, B => n4611, Z => n4934);
   U4590 : AO7 port map( A => n4950, B => n4853, C => n4951, Z => n4200);
   U4591 : AO2 port map( A => n4952, B => n4709, C => n7819, D => n4953, Z => 
                           n4951);
   U4592 : AO7 port map( A => n4954, B => n4853, C => n4955, Z => n4199);
   U4593 : AO2 port map( A => n4952, B => n4714, C => n7818, D => n4953, Z => 
                           n4955);
   U4594 : AO7 port map( A => n4956, B => n4853, C => n4957, Z => n4198);
   U4595 : AO2 port map( A => n4952, B => n4717, C => n7817, D => n4953, Z => 
                           n4957);
   U4596 : AO7 port map( A => n4958, B => n4853, C => n4959, Z => n4197);
   U4597 : AO2 port map( A => n4952, B => n4720, C => n7856, D => n4953, Z => 
                           n4959);
   U4598 : AO7 port map( A => n4960, B => n4853, C => n4961, Z => n4196);
   U4599 : AO2 port map( A => n4952, B => n4723, C => n7816, D => n4953, Z => 
                           n4961);
   U4600 : AO7 port map( A => n4962, B => n4853, C => n4963, Z => n4195);
   U4601 : AO2 port map( A => n4964, B => n4952, C => n7869, D => n4953, Z => 
                           n4963);
   U4602 : MUX21L port map( A => n4965, B => n4966, S => n4396, Z => n4964);
   U4603 : AO1 port map( A => n4967, B => n4968, C => n4969, D => n4970, Z => 
                           n4965);
   U4604 : AO4 port map( A => n4971, B => n4972, C => n4973, D => n4974, Z => 
                           n4970);
   U4605 : AO6 port map( A => n4975, B => n4976, C => n4977, Z => n4973);
   U4606 : AO4 port map( A => n4359, B => n4978, C => n4979, D => n4980, Z => 
                           n4977);
   U4607 : AO4 port map( A => n4404, B => n4981, C => n4982, D => n4983, Z => 
                           n4969);
   U4608 : AO7 port map( A => n4984, B => n4853, C => n4985, Z => n4194);
   U4609 : AO2 port map( A => n4952, B => n4729, C => n7860, D => n4953, Z => 
                           n4985);
   U4610 : AO7 port map( A => n4986, B => n4853, C => n4987, Z => n4193);
   U4611 : AO2 port map( A => n4988, B => n4952, C => n7815, D => n4953, Z => 
                           n4987);
   U4612 : NR2 port map( A => n4911, B => n4953, Z => n4952);
   U4613 : NR2 port map( A => n4911, B => n4658, Z => n4953);
   U4614 : MUX21L port map( A => n4989, B => n4990, S => n4396, Z => n4988);
   U4615 : NR2 port map( A => n4991, B => n4992, Z => n4990);
   U4616 : AN3 port map( A => n4993, B => n4994, C => n4995, Z => n4991);
   U4617 : MUX21L port map( A => n4996, B => n4997, S => n4359, Z => n4995);
   U4618 : AO6 port map( A => n4998, B => v_RAM_OUT0_29_port, C => n4999, Z => 
                           n4989);
   U4619 : AO4 port map( A => n4974, B => n5000, C => n4982, D => n5001, Z => 
                           n4999);
   U4620 : MUX21L port map( A => n5002, B => n5003, S => n5004, Z => n5001);
   U4621 : MUX21L port map( A => n5005, B => n5006, S => n4359, Z => n5002);
   U4622 : IV port map( A => n5007, Z => n4998);
   U4623 : IV port map( A => n4911, Z => n4853);
   U4624 : AO7 port map( A => n5008, B => n5009, C => n5010, Z => n4192);
   U4625 : AO2 port map( A => n5011, B => n4586, C => n7902, D => n5012, Z => 
                           n5010);
   U4626 : IV port map( A => n5013, Z => n4586);
   U4627 : AO7 port map( A => n5014, B => n5015, C => n5016, Z => n5013);
   U4628 : MUX21L port map( A => n5017, B => n5018, S => n4394, Z => n5016);
   U4629 : AO3 port map( A => n4900, B => n5019, C => n5020, D => n5021, Z => 
                           n5018);
   U4630 : AO1 port map( A => n5022, B => n5023, C => n5024, D => n5025, Z => 
                           n5021);
   U4631 : AO6 port map( A => n5026, B => n5027, C => n5028, Z => n5025);
   U4632 : ND3 port map( A => v_RAM_OUT0_2_port, B => n4878, C => n5029, Z => 
                           n5027);
   U4633 : AN3 port map( A => n5030, B => n4360, C => n4873, Z => n5024);
   U4634 : EO1 port map( A => n4907, B => n5031, C => n4870, D => n5032, Z => 
                           n5020);
   U4635 : NR4 port map( A => n5033, B => n5034, C => n5035, D => n5036, Z => 
                           n5017);
   U4636 : AO4 port map( A => n5037, B => n5038, C => n4870, D => n5039, Z => 
                           n5036);
   U4637 : ND2 port map( A => n4887, B => n5040, Z => n5039);
   U4638 : ND2 port map( A => n5041, B => n4406, Z => n5038);
   U4639 : AN3 port map( A => n5042, B => n5043, C => n5044, Z => n5035);
   U4640 : AO4 port map( A => n5045, B => n5046, C => n5047, D => n5048, Z => 
                           n5034);
   U4641 : AO1 port map( A => n5049, B => n4873, C => n5050, D => n5051, Z => 
                           n5045);
   U4642 : AO6 port map( A => n5052, B => n5053, C => n5037, Z => n5051);
   U4643 : AO4 port map( A => n5028, B => n5054, C => n5032, D => n5055, Z => 
                           n5050);
   U4644 : NR2 port map( A => n5056, B => n5057, Z => n5032);
   U4645 : AO3 port map( A => n5058, B => n5026, C => n5059, D => n5060, Z => 
                           n5033);
   U4646 : AO2 port map( A => n5061, B => n5062, C => n5063, D => n5064, Z => 
                           n5060);
   U4647 : AO3 port map( A => n5054, B => n5065, C => n5066, D => n5067, Z => 
                           n5064);
   U4648 : ND2 port map( A => n5068, B => n5069, Z => n5067);
   U4649 : OR3 port map( A => n5070, B => n5071, C => n5055, Z => n5066);
   U4650 : AO4 port map( A => n5055, B => n5072, C => n5073, D => n5037, Z => 
                           n5062);
   U4651 : MUX21L port map( A => n4907, B => n5074, S => n5075, Z => n5059);
   U4652 : NR4 port map( A => n5076, B => n5077, C => n5078, D => n5079, Z => 
                           n5014);
   U4653 : AO4 port map( A => n5080, B => n4897, C => n5081, D => n5040, Z => 
                           n5079);
   U4654 : AO4 port map( A => n5082, B => n5083, C => n5084, D => n5085, Z => 
                           n5078);
   U4655 : AO4 port map( A => n5086, B => n5087, C => n4360, D => n5088, Z => 
                           n5077);
   U4656 : MUX21L port map( A => n4896, B => n5089, S => n4362, Z => n5088);
   U4657 : AO4 port map( A => n5090, B => n5091, C => n4898, D => n5092, Z => 
                           n5076);
   U4658 : OR2 port map( A => n5093, B => n5094, Z => n5092);
   U4659 : AO7 port map( A => n5095, B => n5009, C => n5096, Z => n4191);
   U4660 : AO2 port map( A => n5011, B => n4591, C => n7908, D => n5012, Z => 
                           n5096);
   U4661 : MUX21L port map( A => n5097, B => n5098, S => n4394, Z => n4591);
   U4662 : AO1 port map( A => n5099, B => n5100, C => n5101, D => n5102, Z => 
                           n5098);
   U4663 : AO1 port map( A => n5044, B => n5103, C => n5104, D => n5105, Z => 
                           n5102);
   U4664 : AO4 port map( A => n5106, B => n5107, C => n5108, D => n4880, Z => 
                           n5105);
   U4665 : NR2 port map( A => n5073, B => n5089, Z => n5108);
   U4666 : AO7 port map( A => n5109, B => n5046, C => n4878, Z => n5104);
   U4667 : AO4 port map( A => n5110, B => n5037, C => n5111, D => n5055, Z => 
                           n5101);
   U4668 : AO1 port map( A => n4885, B => n4899, C => n5112, D => n5113, Z => 
                           n5111);
   U4669 : NR2 port map( A => v_RAM_OUT0_4_port, B => n5023, Z => n5113);
   U4670 : AO3 port map( A => n5114, B => n5115, C => n5116, D => n5117, Z => 
                           n5112);
   U4671 : AN3 port map( A => n5118, B => n5119, C => n5063, Z => n5116);
   U4672 : AO1 port map( A => n5120, B => n5061, C => n5121, D => n5122, Z => 
                           n5110);
   U4673 : AO4 port map( A => n5115, B => n5123, C => n5124, D => n5046, Z => 
                           n5121);
   U4674 : NR2 port map( A => n5089, B => n4884, Z => n5124);
   U4675 : NR2 port map( A => n5071, B => n5125, Z => n5120);
   U4676 : AO1 port map( A => n5125, B => n5063, C => n5126, D => n5127, Z => 
                           n5100);
   U4677 : NR2 port map( A => n5046, B => n5128, Z => n5127);
   U4678 : NR2 port map( A => n5129, B => n5130, Z => n5099);
   U4679 : MUX21L port map( A => n5115, B => n5106, S => n5131, Z => n5130);
   U4680 : MUX21L port map( A => n5132, B => n5133, S => n4402, Z => n5097);
   U4681 : AN3 port map( A => n5134, B => n5135, C => n5136, Z => n5133);
   U4682 : AO1 port map( A => n5137, B => n5138, C => n5139, D => n5140, Z => 
                           n5136);
   U4683 : NR4 port map( A => v_RAM_OUT0_2_port, B => v_RAM_OUT0_1_port, C => 
                           n5109, D => n4896, Z => n5140);
   U4684 : AO4 port map( A => n4898, B => n5141, C => n5085, D => n5142, Z => 
                           n5139);
   U4685 : NR2 port map( A => n5069, B => n5143, Z => n5137);
   U4686 : AO2 port map( A => n5144, B => n5145, C => n5094, D => n5146, Z => 
                           n5135);
   U4687 : EO1 port map( A => n5147, B => n5058, C => n5148, D => n5149, Z => 
                           n5134);
   U4688 : NR4 port map( A => n5150, B => n5151, C => n5152, D => n5153, Z => 
                           n5132);
   U4689 : AO4 port map( A => n5090, B => n5154, C => v_RAM_OUT0_1_port, D => 
                           n5052, Z => n5153);
   U4690 : MUX21L port map( A => n5085, B => n5155, S => n4887, Z => n5152);
   U4691 : AO6 port map( A => n5146, B => n5040, C => n5156, Z => n5155);
   U4692 : AO4 port map( A => n5053, B => n5087, C => n5157, D => n5158, Z => 
                           n5151);
   U4693 : AO6 port map( A => n5159, B => n5160, C => n5138, Z => n5158);
   U4694 : AO6 port map( A => n5019, B => n5123, C => n5081, Z => n5150);
   U4695 : AO7 port map( A => n5161, B => n5009, C => n5162, Z => n4190);
   U4696 : AO2 port map( A => n5011, B => n4594, C => n7914, D => n5012, Z => 
                           n5162);
   U4697 : MUX21H port map( A => n5163, B => n5164, S => v_RAM_OUT0_7_port, Z 
                           => n4594);
   U4698 : AO1 port map( A => n5165, B => n5166, C => n5167, D => n5168, Z => 
                           n5164);
   U4699 : AO4 port map( A => n5040, B => n4900, C => n5169, D => n5055, Z => 
                           n5168);
   U4700 : AO1 port map( A => n4885, B => n4908, C => n5170, D => n5171, Z => 
                           n5169);
   U4701 : AO7 port map( A => n5106, B => n5172, C => n5173, Z => n5171);
   U4702 : IV port map( A => n5122, Z => n5173);
   U4703 : AO4 port map( A => n5115, B => n5174, C => n4880, D => n4886, Z => 
                           n5170);
   U4704 : AO3 port map( A => n5175, B => n5037, C => n5176, D => n5177, Z => 
                           n5167);
   U4705 : AO2 port map( A => n5178, B => n5179, C => n5180, D => n4873, Z => 
                           n5177);
   U4706 : AO7 port map( A => n4907, B => n5074, C => n4884, Z => n5176);
   U4707 : AO1 port map( A => n5061, B => n4908, C => n5181, D => n5182, Z => 
                           n5175);
   U4708 : IV port map( A => n5183, Z => n5182);
   U4709 : AO6 port map( A => n5184, B => n5044, C => n5185, Z => n5183);
   U4710 : AO4 port map( A => n4880, B => n5031, C => n5046, D => n5072, Z => 
                           n5181);
   U4711 : AO1 port map( A => n5061, B => n5186, C => n5185, D => n5187, Z => 
                           n5166);
   U4712 : AO6 port map( A => n5119, B => n5188, C => n5046, Z => n5187);
   U4713 : ND2 port map( A => n5023, B => n5189, Z => n5186);
   U4714 : AO1 port map( A => n5044, B => n5190, C => n5054, D => n5191, Z => 
                           n5165);
   U4715 : NR2 port map( A => n4880, B => n5192, Z => n5191);
   U4716 : AO7 port map( A => n5193, B => n5037, C => n5194, Z => n5163);
   U4717 : MUX21L port map( A => n5195, B => n5196, S => n4402, Z => n5194);
   U4718 : NR4 port map( A => n5197, B => n5198, C => n5199, D => n5200, Z => 
                           n5196);
   U4719 : AO4 port map( A => n5082, B => n5081, C => n5072, D => n5149, Z => 
                           n5200);
   U4720 : MUX21L port map( A => n4897, B => n5087, S => n4908, Z => n5199);
   U4721 : AO4 port map( A => n5090, B => n5201, C => n5202, D => n4898, Z => 
                           n5198);
   U4722 : IV port map( A => n5203, Z => n4898);
   U4723 : ND2 port map( A => n5204, B => n5019, Z => n5201);
   U4724 : EON1 port map( A => n5205, B => n5085, C => n5206, D => n5159, Z => 
                           n5197);
   U4725 : AO4 port map( A => n5207, B => n5208, C => n5081, D => n5192, Z => 
                           n5195);
   U4726 : AO7 port map( A => n5209, B => n5106, C => n5210, Z => n5208);
   U4727 : AO3 port map( A => n5049, B => n5115, C => n4883, D => n4362, Z => 
                           n5207);
   U4728 : IV port map( A => n5126, Z => n4883);
   U4729 : NR2 port map( A => n5211, B => n5046, Z => n5126);
   U4730 : AO1 port map( A => n5212, B => n5063, C => n5213, D => n5214, Z => 
                           n5193);
   U4731 : NR3 port map( A => n5115, B => n4896, C => n5093, Z => n5214);
   U4732 : NR2 port map( A => n4360, B => n5119, Z => n5213);
   U4733 : AO7 port map( A => n5215, B => n5009, C => n5216, Z => n4189);
   U4734 : AO2 port map( A => n5011, B => n4597, C => n7920, D => n5012, Z => 
                           n5216);
   U4735 : MUX21L port map( A => n5217, B => n5218, S => n4394, Z => n4597);
   U4736 : AO1 port map( A => n5219, B => n5220, C => n5221, D => n5222, Z => 
                           n5218);
   U4737 : AO1 port map( A => n5084, B => n5063, C => n5223, D => n5224, Z => 
                           n5222);
   U4738 : AO4 port map( A => n5115, B => n5192, C => n5225, D => n5046, Z => 
                           n5224);
   U4739 : AO7 port map( A => n5106, B => n4908, C => n4878, Z => n5223);
   U4740 : AO4 port map( A => n5226, B => n5055, C => n5227, D => n5037, Z => 
                           n5221);
   U4741 : AO1 port map( A => n5061, B => n5228, C => n5229, D => n5230, Z => 
                           n5227);
   U4742 : AN3 port map( A => n4885, B => n5075, C => n5231, Z => n5230);
   U4743 : AO4 port map( A => n4880, B => n5211, C => n5115, D => n4901, Z => 
                           n5229);
   U4744 : ND2 port map( A => n5031, B => n5052, Z => n5228);
   U4745 : AO1 port map( A => n5061, B => n5107, C => n5232, D => n5233, Z => 
                           n5226);
   U4746 : AO6 port map( A => n5231, B => n5019, C => n5115, Z => n5233);
   U4747 : AO4 port map( A => n5046, B => n5118, C => n4880, D => n5047, Z => 
                           n5232);
   U4748 : IV port map( A => n5234, Z => n5107);
   U4749 : AO1 port map( A => n4885, B => n5235, C => n5185, D => n5122, Z => 
                           n5220);
   U4750 : NR2 port map( A => n5023, B => n4880, Z => n5122);
   U4751 : NR2 port map( A => n5072, B => n4880, Z => n5185);
   U4752 : AO1 port map( A => n5202, B => n5061, C => n5129, D => n5236, Z => 
                           n5219);
   U4753 : AO6 port map( A => n5237, B => n5043, C => n5115, Z => n5236);
   U4754 : AO1 port map( A => n5068, B => n5238, C => n5239, D => n5240, Z => 
                           n5217);
   U4755 : AO4 port map( A => n5241, B => n5055, C => n5242, D => n5054, Z => 
                           n5240);
   U4756 : AO1 port map( A => n5184, B => n4360, C => n5243, D => n5244, Z => 
                           n5242);
   U4757 : AN3 port map( A => n5128, B => n5119, C => n4885, Z => n5244);
   U4758 : NR2 port map( A => v_RAM_OUT0_4_port, B => n5131, Z => n5243);
   U4759 : IV port map( A => n5042, Z => n5055);
   U4760 : AO1 port map( A => n5061, B => n5142, C => n5245, D => n5180, Z => 
                           n5241);
   U4761 : NR2 port map( A => n5142, B => n5046, Z => n5180);
   U4762 : AO4 port map( A => n4880, B => n5204, C => v_RAM_OUT0_2_port, D => 
                           n5023, Z => n5245);
   U4763 : IV port map( A => n5246, Z => n5142);
   U4764 : ND4 port map( A => n5247, B => n5248, C => n5249, D => n4870, Z => 
                           n5239);
   U4765 : ND4 port map( A => n5044, B => n4886, C => n5023, D => n4402, Z => 
                           n5249);
   U4766 : IV port map( A => n5057, Z => n5023);
   U4767 : OR3 port map( A => n5029, B => n5250, C => n4900, Z => n5248);
   U4768 : AO7 port map( A => n5251, B => n4907, C => n5188, Z => n5247);
   U4769 : AN3 port map( A => n4873, B => v_RAM_OUT0_4_port, C => n5093, Z => 
                           n5251);
   U4770 : AO3 port map( A => n5106, B => n5252, C => n5253, D => n5254, Z => 
                           n5238);
   U4771 : AO2 port map( A => n5063, B => n5255, C => n5256, D => n5044, Z => 
                           n5254);
   U4772 : ND2 port map( A => n5174, B => n5145, Z => n5255);
   U4773 : ND3 port map( A => n5123, B => n5019, C => n4885, Z => n5253);
   U4774 : ND2 port map( A => n5128, B => n5119, Z => n5252);
   U4775 : AO7 port map( A => n5257, B => n5009, C => n5258, Z => n4188);
   U4776 : AO2 port map( A => n5011, B => n4600, C => n7926, D => n5012, Z => 
                           n5258);
   U4777 : IV port map( A => n5259, Z => n4600);
   U4778 : AO7 port map( A => n5260, B => n5015, C => n5261, Z => n5259);
   U4779 : MUX21L port map( A => n5262, B => n5263, S => n4394, Z => n5261);
   U4780 : ND4 port map( A => n5264, B => n5265, C => n5266, D => n5267, Z => 
                           n5263);
   U4781 : AO2 port map( A => n4876, B => n5268, C => n5269, D => n5270, Z => 
                           n5267);
   U4782 : ND2 port map( A => n5204, B => n5192, Z => n5268);
   U4783 : IV port map( A => n5271, Z => n5266);
   U4784 : AO4 port map( A => n5272, B => n5128, C => n5141, D => n5273, Z => 
                           n5271);
   U4785 : AO2 port map( A => n5178, B => n5172, C => n4907, D => n5040, Z => 
                           n5265);
   U4786 : ND2 port map( A => n5019, B => n4886, Z => n5172);
   U4787 : IV port map( A => n5080, Z => n4886);
   U4788 : IV port map( A => n5274, Z => n5264);
   U4789 : AO4 port map( A => n4870, B => n5157, C => n4900, D => n5084, Z => 
                           n5274);
   U4790 : NR2 port map( A => n5160, B => n5073, Z => n5157);
   U4791 : NR4 port map( A => n5275, B => n5276, C => n5277, D => n5278, Z => 
                           n5262);
   U4792 : AO4 port map( A => n5279, B => n5280, C => n5109, D => n4900, Z => 
                           n5278);
   U4793 : AO3 port map( A => n5281, B => n5149, C => v_RAM_OUT0_5_port, D => 
                           n5282, Z => n5280);
   U4794 : EO1 port map( A => n5283, B => n5047, C => n5087, D => n5284, Z => 
                           n5282);
   U4795 : IV port map( A => n5028, Z => n5047);
   U4796 : NR2 port map( A => n4881, B => n5071, Z => n5028);
   U4797 : AO3 port map( A => n5285, B => n5090, C => n5286, D => n5287, Z => 
                           n5279);
   U4798 : AO2 port map( A => n5147, B => n5288, C => n5146, D => n5289, Z => 
                           n5287);
   U4799 : ND2 port map( A => n5237, B => n5040, Z => n5289);
   U4800 : ND2 port map( A => n5188, B => n5179, Z => n5288);
   U4801 : AO2 port map( A => n5290, B => n5138, C => n5291, D => n5203, Z => 
                           n5286);
   U4802 : NR2 port map( A => n4896, B => n5160, Z => n5290);
   U4803 : NR2 port map( A => n5029, B => n5292, Z => n5285);
   U4804 : AO4 port map( A => n5040, B => n5026, C => n5293, D => n5148, Z => 
                           n5277);
   U4805 : AO4 port map( A => n5048, B => n5058, C => n5273, D => n5294, Z => 
                           n5276);
   U4806 : AO3 port map( A => n5125, B => n5272, C => n5295, D => n5296, Z => 
                           n5275);
   U4807 : ND3 port map( A => n5174, B => n5145, C => n5270, Z => n5296);
   U4808 : OR3 port map( A => n5269, B => n5143, C => n4870, Z => n5295);
   U4809 : AO1 port map( A => n5297, B => n5188, C => n5298, D => n5299, Z => 
                           n5260);
   U4810 : AO4 port map( A => n5300, B => n5301, C => n5081, D => n5091, Z => 
                           n5299);
   U4811 : ND2 port map( A => n5211, B => n4887, Z => n5091);
   U4812 : IV port map( A => n4884, Z => n4887);
   U4813 : AO6 port map( A => n5159, B => n5302, C => n5138, Z => n5300);
   U4814 : NR2 port map( A => n4362, B => v_RAM_OUT0_2_port, Z => n5159);
   U4815 : AO7 port map( A => n5281, B => n5085, C => n5303, Z => n5298);
   U4816 : AO2 port map( A => n5156, B => n5302, C => n5250, D => n5304, Z => 
                           n5303);
   U4817 : ND2 port map( A => n5128, B => n5043, Z => n5302);
   U4818 : AO7 port map( A => n5069, B => n5087, C => n4897, Z => n5297);
   U4819 : AO7 port map( A => n5305, B => n5009, C => n5306, Z => n4187);
   U4820 : AO2 port map( A => n5307, B => n5011, C => n7932, D => n5012, Z => 
                           n5306);
   U4821 : MUX21L port map( A => n5308, B => n4868, S => n4394, Z => n5307);
   U4822 : ND4 port map( A => n5309, B => n5310, C => n5311, D => n5312, Z => 
                           n4868);
   U4823 : AO1 port map( A => n5042, B => n5313, C => n5314, D => n5315, Z => 
                           n5312);
   U4824 : AO4 port map( A => n5316, B => n5037, C => n5284, D => n4870, Z => 
                           n5315);
   U4825 : NR2 port map( A => n5317, B => n5056, Z => n5284);
   U4826 : IV port map( A => n5068, Z => n5037);
   U4827 : NR2 port map( A => n5318, B => n5319, Z => n5316);
   U4828 : AO4 port map( A => n5205, B => n4880, C => n5106, D => n5206, Z => 
                           n5319);
   U4829 : ND2 port map( A => n5281, B => n5192, Z => n5206);
   U4830 : EON1 port map( A => n5225, B => n5046, C => n5320, D => n5044, Z => 
                           n5318);
   U4831 : NR2 port map( A => n5071, B => n5269, Z => n5225);
   U4832 : AO4 port map( A => n5026, B => n5145, C => n5293, D => n5204, Z => 
                           n5314);
   U4833 : IV port map( A => n5321, Z => n5145);
   U4834 : AO3 port map( A => n5046, B => n5231, C => n5210, D => n5322, Z => 
                           n5313);
   U4835 : AO2 port map( A => n5044, B => n5323, C => n5061, D => n5324, Z => 
                           n5322);
   U4836 : ND2 port map( A => n5192, B => n5189, Z => n5324);
   U4837 : ND2 port map( A => n5019, B => n5052, Z => n5323);
   U4838 : IV port map( A => n5114, Z => n5052);
   U4839 : AO2 port map( A => n4885, B => n5143, C => n5141, D => n5063, Z => 
                           n5210);
   U4840 : ND2 port map( A => n5231, B => n5053, Z => n5141);
   U4841 : AO2 port map( A => n5270, B => n5202, C => n5325, D => n5109, Z => 
                           n5311);
   U4842 : AO7 port map( A => n5022, B => n4907, C => n5326, Z => n5310);
   U4843 : AO2 port map( A => n5327, B => n5074, C => n5328, D => n5329, Z => 
                           n5309);
   U4844 : ND2 port map( A => n5026, B => n5048, Z => n5329);
   U4845 : NR2 port map( A => n5094, B => n5093, Z => n5327);
   U4846 : AO1 port map( A => n5330, B => n4876, C => n5331, D => n5332, Z => 
                           n5308);
   U4847 : AO4 port map( A => n4870, B => n5154, C => n5333, D => n5054, Z => 
                           n5332);
   U4848 : AO6 port map( A => n5317, B => v_RAM_OUT0_2_port, C => n5334, Z => 
                           n5333);
   U4849 : AO4 port map( A => n5109, B => n4880, C => n5046, D => n5043, Z => 
                           n5334);
   U4850 : AO4 port map( A => n4402, B => n4875, C => n5129, D => n4874, Z => 
                           n5331);
   U4851 : AO3 port map( A => n5335, B => n5188, C => n5336, D => n5337, Z => 
                           n4874);
   U4852 : AO2 port map( A => n5114, B => n4885, C => n5041, D => n5063, Z => 
                           n5337);
   U4853 : NR2 port map( A => n5179, B => v_RAM_OUT0_0_port, Z => n5114);
   U4854 : ND2 port map( A => n5044, B => n5131, Z => n5336);
   U4855 : ND4 port map( A => n5338, B => n5339, C => n5340, D => n5341, Z => 
                           n4875);
   U4856 : AO2 port map( A => n5342, B => n5283, C => n5304, D => n5343, Z => 
                           n5341);
   U4857 : ND2 port map( A => n5075, B => n5189, Z => n5343);
   U4858 : IV port map( A => n5269, Z => n5189);
   U4859 : NR2 port map( A => n4365, B => v_RAM_OUT0_0_port, Z => n5269);
   U4860 : NR2 port map( A => n5321, B => n5330, Z => n5342);
   U4861 : AO2 port map( A => n5203, B => n5103, C => n5144, D => n5344, Z => 
                           n5340);
   U4862 : ND2 port map( A => n5128, B => n5117, Z => n5103);
   U4863 : AO2 port map( A => n5138, B => n5075, C => n5147, D => n5148, Z => 
                           n5339);
   U4864 : AO2 port map( A => n5146, B => n5204, C => n5156, D => n5040, Z => 
                           n5338);
   U4865 : AO7 port map( A => n5345, B => n5009, C => n5346, Z => n4186);
   U4866 : AO2 port map( A => n5011, B => n4606, C => n7938, D => n5012, Z => 
                           n5346);
   U4867 : IV port map( A => n5347, Z => n4606);
   U4868 : AO7 port map( A => n5348, B => n5015, C => n5349, Z => n5347);
   U4869 : MUX21L port map( A => n5350, B => n5351, S => n4394, Z => n5349);
   U4870 : ND4 port map( A => n5352, B => n5353, C => n5354, D => n5355, Z => 
                           n5351);
   U4871 : AO2 port map( A => n5291, B => n5325, C => n5178, D => n5356, Z => 
                           n5355);
   U4872 : ND2 port map( A => n5118, B => n5281, Z => n5356);
   U4873 : NR2 port map( A => n5125, B => n5317, Z => n5291);
   U4874 : AO2 port map( A => n5074, B => n5357, C => n5270, D => n5358, Z => 
                           n5354);
   U4875 : NR2 port map( A => n5054, B => n5046, Z => n5270);
   U4876 : ND2 port map( A => n5031, B => n5040, Z => n5357);
   U4877 : IV port map( A => n5056, Z => n5040);
   U4878 : EO1 port map( A => n5022, B => n5294, C => n5293, D => n5049, Z => 
                           n5353);
   U4879 : NR2 port map( A => n5056, B => n5321, Z => n5049);
   U4880 : ND2 port map( A => n5237, B => n5204, Z => n5294);
   U4881 : IV port map( A => n5359, Z => n5237);
   U4882 : IV port map( A => n5360, Z => n5352);
   U4883 : AO4 port map( A => n4870, B => n5082, C => n5026, D => n5084, Z => 
                           n5360);
   U4884 : IV port map( A => n4876, Z => n5026);
   U4885 : NR4 port map( A => n5361, B => n5362, C => n5363, D => n5364, Z => 
                           n5350);
   U4886 : AO4 port map( A => n5365, B => n5366, C => n5293, D => n5184, Z => 
                           n5364);
   U4887 : OR2 port map( A => n5202, B => n5321, Z => n5184);
   U4888 : IV port map( A => n4907, Z => n5293);
   U4889 : NR2 port map( A => n5129, B => n4880, Z => n4907);
   U4890 : AO3 port map( A => n5069, B => n4897, C => v_RAM_OUT0_5_port, D => 
                           n5367, Z => n5366);
   U4891 : AO2 port map( A => n5147, B => n5154, C => n5205, D => n5144, Z => 
                           n5367);
   U4892 : IV port map( A => n4869, Z => n5154);
   U4893 : NR2 port map( A => n4881, B => n5143, Z => n4869);
   U4894 : AO3 port map( A => n5083, B => n5118, C => n5368, D => n5369, Z => 
                           n5365);
   U4895 : AO2 port map( A => n5250, B => n5203, C => n5283, D => 
                           v_RAM_OUT0_3_port, Z => n5369);
   U4896 : EO1 port map( A => n5370, B => n5304, C => n5149, D => n5086, Z => 
                           n5368);
   U4897 : NR2 port map( A => n5057, B => n5202, Z => n5086);
   U4898 : IV port map( A => n5156, Z => n5149);
   U4899 : NR2 port map( A => n5109, B => n5317, Z => n5370);
   U4900 : MUX21L port map( A => n5272, B => n5371, S => n5058, Z => n5363);
   U4901 : NR2 port map( A => n5372, B => n4876, Z => n5371);
   U4902 : NR2 port map( A => n5054, B => n5106, Z => n4876);
   U4903 : OR3 port map( A => n5330, B => v_RAM_OUT0_2_port, C => n4878, Z => 
                           n5372);
   U4904 : IV port map( A => n5325, Z => n5272);
   U4905 : NR2 port map( A => n5129, B => n5046, Z => n5325);
   U4906 : AO4 port map( A => n4900, B => n5030, C => n5256, D => n5048, Z => 
                           n5362);
   U4907 : IV port map( A => n5178, Z => n5048);
   U4908 : NR2 port map( A => n5129, B => n5115, Z => n5178);
   U4909 : NR2 port map( A => n5069, B => n5321, Z => n5256);
   U4910 : NR2 port map( A => n4881, B => n4356, Z => n5321);
   U4911 : ND2 port map( A => n5174, B => n5373, Z => n5030);
   U4912 : IV port map( A => n5074, Z => n4900);
   U4913 : NR2 port map( A => n5129, B => n5106, Z => n5074);
   U4914 : AO4 port map( A => n5273, B => n5043, C => n4870, D => n5374, Z => 
                           n5361);
   U4915 : ND2 port map( A => n5019, B => n5123, Z => n5374);
   U4916 : IV port map( A => n5041, Z => n5123);
   U4917 : IV port map( A => n5326, Z => n5019);
   U4918 : ND2 port map( A => n4878, B => n5044, Z => n4870);
   U4919 : IV port map( A => n5022, Z => n5273);
   U4920 : NR2 port map( A => n5054, B => n4880, Z => n5022);
   U4921 : ND2 port map( A => v_RAM_OUT0_5_port, B => n4394, Z => n5015);
   U4922 : NR4 port map( A => n5375, B => n5376, C => n5377, D => n5378, Z => 
                           n5348);
   U4923 : AO4 port map( A => n5085, B => n4901, C => n5084, D => n5083, Z => 
                           n5378);
   U4924 : NR2 port map( A => n5359, B => n5093, Z => n5084);
   U4925 : NR2 port map( A => v_RAM_OUT0_0_port, B => n5070, Z => n5093);
   U4926 : IV port map( A => n5212, Z => n4901);
   U4927 : IV port map( A => n5283, Z => n5085);
   U4928 : EON1 port map( A => n5081, B => n5344, C => n5065, D => n5156, Z => 
                           n5377);
   U4929 : IV port map( A => n5147, Z => n5081);
   U4930 : EON1 port map( A => n5379, B => n4897, C => n5190, D => n5203, Z => 
                           n5376);
   U4931 : ND2 port map( A => n5174, B => n5053, Z => n5190);
   U4932 : IV port map( A => n5330, Z => n5174);
   U4933 : IV port map( A => n5146, Z => n4897);
   U4934 : NR2 port map( A => n5041, B => n5029, Z => n5379);
   U4935 : NR2 port map( A => n5281, B => v_RAM_OUT0_0_port, Z => n5041);
   U4936 : AO4 port map( A => n5380, B => n5087, C => n5090, D => n5235, Z => 
                           n5375);
   U4937 : ND2 port map( A => n5192, B => n5131, Z => n5235);
   U4938 : IV port map( A => n5143, Z => n5192);
   U4939 : NR2 port map( A => n4356, B => n5070, Z => n5143);
   U4940 : IV port map( A => n5304, Z => n5090);
   U4941 : IV port map( A => n5144, Z => n5087);
   U4942 : NR2 port map( A => n5056, B => n4896, Z => n5380);
   U4943 : AO7 port map( A => n5381, B => n5009, C => n5382, Z => n4185);
   U4944 : AO2 port map( A => n5383, B => n5011, C => n7944, D => n5012, Z => 
                           n5382);
   U4945 : NR2 port map( A => n5384, B => n5012, Z => n5011);
   U4946 : NR2 port map( A => n5384, B => n4658, Z => n5012);
   U4947 : NR2 port map( A => n5385, B => n4536, Z => n4658);
   U4948 : MUX21L port map( A => n5386, B => n5387, S => n4394, Z => n5383);
   U4949 : NR2 port map( A => n5388, B => n4895, Z => n5387);
   U4950 : AO3 port map( A => n5058, B => n5389, C => n5390, D => n5391, Z => 
                           n4895);
   U4951 : ND4 port map( A => n5392, B => n5393, C => n5394, D => n5395, Z => 
                           n5391);
   U4952 : NR2 port map( A => v_RAM_OUT0_5_port, B => n5396, Z => n5395);
   U4953 : AO6 port map( A => n5075, B => n5231, C => n5115, Z => n5396);
   U4954 : IV port map( A => n5160, Z => n5231);
   U4955 : NR2 port map( A => v_RAM_OUT0_0_port, B => n5069, Z => n5160);
   U4956 : IV port map( A => n4896, Z => n5075);
   U4957 : AO2 port map( A => n5203, B => n5320, C => n5146, D => n5344, Z => 
                           n5394);
   U4958 : ND2 port map( A => n5118, B => n5211, Z => n5344);
   U4959 : IV port map( A => n5071, Z => n5118);
   U4960 : NR2 port map( A => n4356, B => n5069, Z => n5071);
   U4961 : NR2 port map( A => n5106, B => n4362, Z => n5146);
   U4962 : ND2 port map( A => n5211, B => n5188, Z => n5320);
   U4963 : IV port map( A => n5317, Z => n5188);
   U4964 : AO2 port map( A => n5304, B => n5128, C => n5283, D => n5069, Z => 
                           n5393);
   U4965 : AO2 port map( A => n5359, B => n5147, C => n5156, D => n4365, Z => 
                           n5392);
   U4966 : NR2 port map( A => n4356, B => n4407, Z => n5359);
   U4967 : ND3 port map( A => n5042, B => n5397, C => n5398, Z => n5390);
   U4968 : AO1 port map( A => n4896, B => n5044, C => n5056, D => n5399, Z => 
                           n5398);
   U4969 : NR2 port map( A => n4884, B => n5106, Z => n5399);
   U4970 : NR2 port map( A => n5281, B => n4356, Z => n4884);
   U4971 : IV port map( A => n5400, Z => n5281);
   U4972 : NR2 port map( A => v_RAM_OUT0_3_port, B => v_RAM_OUT0_0_port, Z => 
                           n5056);
   U4973 : AO4 port map( A => n5326, B => n5082, C => n5063, D => n5401, Z => 
                           n5397);
   U4974 : NR2 port map( A => v_RAM_OUT0_4_port, B => n5204, Z => n5401);
   U4975 : IV port map( A => n5082, Z => n5204);
   U4976 : NR2 port map( A => v_RAM_OUT0_0_port, B => n5400, Z => n5082);
   U4977 : NR2 port map( A => n4402, B => v_RAM_OUT0_1_port, Z => n5042);
   U4978 : ND2 port map( A => n5068, B => n5335, Z => n5389);
   U4979 : IV port map( A => n5402, Z => n5058);
   U4980 : AN3 port map( A => n4910, B => n5068, C => n5403, Z => n5388);
   U4981 : MUX21L port map( A => n4896, B => n4899, S => n4360, Z => n5403);
   U4982 : IV port map( A => n5209, Z => n4899);
   U4983 : NR2 port map( A => n5029, B => n5080, Z => n5209);
   U4984 : NR2 port map( A => n4881, B => v_RAM_OUT0_0_port, Z => n5080);
   U4985 : NR2 port map( A => n4362, B => n4402, Z => n5068);
   U4986 : AO6 port map( A => n5404, B => v_RAM_OUT0_5_port, C => n5405, Z => 
                           n5386);
   U4987 : AO4 port map( A => n5054, B => n4904, C => n5129, D => n5406, Z => 
                           n5405);
   U4988 : MUX21L port map( A => n5407, B => n4909, S => n5335, Z => n5406);
   U4989 : IV port map( A => n4910, Z => n5335);
   U4990 : NR2 port map( A => n5044, B => n4885, Z => n4910);
   U4991 : IV port map( A => n5301, Z => n4909);
   U4992 : ND2 port map( A => n5211, B => n5053, Z => n5301);
   U4993 : ND2 port map( A => n5069, B => v_RAM_OUT0_0_port, Z => n5053);
   U4994 : MUX21L port map( A => n5212, B => n4908, S => n4360, Z => n5407);
   U4995 : IV port map( A => n5358, Z => n4908);
   U4996 : NR2 port map( A => n5330, B => n5057, Z => n5358);
   U4997 : NR2 port map( A => n4356, B => v_RAM_OUT0_6_port, Z => n5057);
   U4998 : NR2 port map( A => n4896, B => n5070, Z => n5212);
   U4999 : IV port map( A => n4873, Z => n5129);
   U5000 : NR2 port map( A => n4362, B => v_RAM_OUT0_5_port, Z => n4873);
   U5001 : AO7 port map( A => n5246, B => n5115, C => n5408, Z => n4904);
   U5002 : AO2 port map( A => n5402, B => n5409, C => n5234, D => n5063, Z => 
                           n5408);
   U5003 : AO7 port map( A => n4360, B => n5117, C => n5106, Z => n5409);
   U5004 : IV port map( A => n5089, Z => n5117);
   U5005 : NR2 port map( A => n5326, B => n5330, Z => n5402);
   U5006 : NR2 port map( A => v_RAM_OUT0_0_port, B => n5109, Z => n5330);
   U5007 : NR2 port map( A => n4356, B => v_RAM_OUT0_3_port, Z => n5326);
   U5008 : NR2 port map( A => n5073, B => n5202, Z => n5246);
   U5009 : NR2 port map( A => n5119, B => v_RAM_OUT0_0_port, Z => n5202);
   U5010 : IV port map( A => n4878, Z => n5054);
   U5011 : NR2 port map( A => v_RAM_OUT0_5_port, B => v_RAM_OUT0_1_port, Z => 
                           n4878);
   U5012 : IV port map( A => n4905, Z => n5404);
   U5013 : ND4 port map( A => n5410, B => n5411, C => n5412, D => n5413, Z => 
                           n4905);
   U5014 : AO2 port map( A => v_RAM_OUT0_1_port, B => n5414, C => n5234, D => 
                           n5283, Z => n5413);
   U5015 : NR2 port map( A => n5046, B => v_RAM_OUT0_1_port, Z => n5283);
   U5016 : NR2 port map( A => n4896, B => n5400, Z => n5234);
   U5017 : NR2 port map( A => n4356, B => n5125, Z => n4896);
   U5018 : AO4 port map( A => n4406, B => n5072, C => n5415, D => n4360, Z => 
                           n5414);
   U5019 : NR2 port map( A => n5089, B => n5094, Z => n5415);
   U5020 : NR2 port map( A => n5131, B => v_RAM_OUT0_0_port, Z => n5089);
   U5021 : IV port map( A => n5069, Z => n5131);
   U5022 : NR2 port map( A => n4365, B => v_RAM_OUT0_6_port, Z => n5069);
   U5023 : IV port map( A => n5250, Z => n5072);
   U5024 : NR2 port map( A => v_RAM_OUT0_0_port, B => n5125, Z => n5250);
   U5025 : EO1 port map( A => n5144, B => n5065, C => n5083, D => n5205, Z => 
                           n5412);
   U5026 : NR2 port map( A => n5073, B => n5328, Z => n5205);
   U5027 : NR2 port map( A => n4365, B => n4356, Z => n5073);
   U5028 : IV port map( A => n5138, Z => n5083);
   U5029 : NR2 port map( A => n5115, B => n4362, Z => n5138);
   U5030 : ND2 port map( A => n5211, B => n5373, Z => n5065);
   U5031 : IV port map( A => n5094, Z => n5373);
   U5032 : NR2 port map( A => n4356, B => n5179, Z => n5094);
   U5033 : IV port map( A => n5070, Z => n5179);
   U5034 : NR2 port map( A => n4407, B => v_RAM_OUT0_3_port, Z => n5070);
   U5035 : IV port map( A => n5292, Z => n5211);
   U5036 : NR2 port map( A => n4407, B => v_RAM_OUT0_0_port, Z => n5292);
   U5037 : NR2 port map( A => n5115, B => v_RAM_OUT0_1_port, Z => n5144);
   U5038 : IV port map( A => n5044, Z => n5115);
   U5039 : NR2 port map( A => v_RAM_OUT0_4_port, B => v_RAM_OUT0_2_port, Z => 
                           n5044);
   U5040 : AO2 port map( A => n5304, B => n5148, C => n5203, D => n5128, Z => 
                           n5411);
   U5041 : ND2 port map( A => v_RAM_OUT0_0_port, B => n4881, Z => n5128);
   U5042 : IV port map( A => n5109, Z => n4881);
   U5043 : NR2 port map( A => n4362, B => n4880, Z => n5203);
   U5044 : ND2 port map( A => n5031, B => n5043, Z => n5148);
   U5045 : IV port map( A => n5328, Z => n5043);
   U5046 : NR2 port map( A => v_RAM_OUT0_6_port, B => v_RAM_OUT0_0_port, Z => 
                           n5328);
   U5047 : IV port map( A => n5029, Z => n5031);
   U5048 : NR2 port map( A => n5119, B => n4356, Z => n5029);
   U5049 : IV port map( A => n5125, Z => n5119);
   U5050 : NR2 port map( A => n4880, B => v_RAM_OUT0_1_port, Z => n5304);
   U5051 : IV port map( A => n5063, Z => n4880);
   U5052 : NR2 port map( A => n4406, B => v_RAM_OUT0_2_port, Z => n5063);
   U5053 : AO2 port map( A => n5156, B => n5109, C => n5317, D => n5147, Z => 
                           n5410);
   U5054 : NR2 port map( A => n5046, B => n4362, Z => n5147);
   U5055 : IV port map( A => n4885, Z => n5046);
   U5056 : NR2 port map( A => n4360, B => n4406, Z => n4885);
   U5057 : NR2 port map( A => n4356, B => n5400, Z => n5317);
   U5058 : NR2 port map( A => n5125, B => n5400, Z => n5109);
   U5059 : NR2 port map( A => n4365, B => n4407, Z => n5400);
   U5060 : NR2 port map( A => v_RAM_OUT0_6_port, B => v_RAM_OUT0_3_port, Z => 
                           n5125);
   U5061 : NR2 port map( A => n5106, B => v_RAM_OUT0_1_port, Z => n5156);
   U5062 : IV port map( A => n5061, Z => n5106);
   U5063 : NR2 port map( A => n4360, B => v_RAM_OUT0_4_port, Z => n5061);
   U5064 : AO7 port map( A => n5416, B => n5009, C => n5417, Z => n4184);
   U5065 : AO2 port map( A => n5418, B => n4615, C => n7814, D => n5419, Z => 
                           n5417);
   U5066 : AO6 port map( A => n5420, B => n5421, C => n5422, Z => n4615);
   U5067 : MUX21H port map( A => n5423, B => n5424, S => v_RAM_OUT0_9_port, Z 
                           => n5422);
   U5068 : NR2 port map( A => v_RAM_OUT0_15_port, B => n5425, Z => n5424);
   U5069 : NR4 port map( A => n5426, B => n5427, C => n5428, D => n5429, Z => 
                           n5425);
   U5070 : AO4 port map( A => n5430, B => n5431, C => n5432, D => n5433, Z => 
                           n5429);
   U5071 : AO4 port map( A => n5434, B => n5435, C => n5436, D => n5437, Z => 
                           n5428);
   U5072 : AO4 port map( A => n5438, B => n4649, C => n5439, D => n5440, Z => 
                           n5427);
   U5073 : NR2 port map( A => n5441, B => n5442, Z => n5439);
   U5074 : AO4 port map( A => n4353, B => n5443, C => n5444, D => n5445, Z => 
                           n5426);
   U5075 : ND2 port map( A => n5446, B => n5447, Z => n5445);
   U5076 : ND2 port map( A => v_RAM_OUT0_8_port, B => n4398, Z => n5443);
   U5077 : AO3 port map( A => n5448, B => n5449, C => n5450, D => n5451, Z => 
                           n5423);
   U5078 : AO2 port map( A => n4665, B => n5452, C => n5453, D => n5454, Z => 
                           n5451);
   U5079 : AO3 port map( A => n5455, B => n5456, C => n5457, D => n5458, Z => 
                           n5454);
   U5080 : AO2 port map( A => n5459, B => v_RAM_OUT0_10_port, C => n5460, D => 
                           n5461, Z => n5458);
   U5081 : OR2 port map( A => n5462, B => n5463, Z => n5457);
   U5082 : AO7 port map( A => n5464, B => n5465, C => n5466, Z => n5452);
   U5083 : AO2 port map( A => n5467, B => n5468, C => n5469, D => n5470, Z => 
                           n5466);
   U5084 : AO7 port map( A => n4357, B => n5471, C => n5432, Z => n5467);
   U5085 : OR3 port map( A => n5472, B => n5464, C => n5470, Z => n5450);
   U5086 : AO3 port map( A => n4676, B => n5473, C => v_RAM_OUT0_15_port, D => 
                           n5474, Z => n5449);
   U5087 : AO2 port map( A => n5475, B => n5476, C => n5477, D => n5478, Z => 
                           n5474);
   U5088 : AO3 port map( A => n5479, B => n5480, C => n5481, D => n5482, Z => 
                           n5448);
   U5089 : AO2 port map( A => n5483, B => n5484, C => n5485, D => n5468, Z => 
                           n5482);
   U5090 : ND2 port map( A => n5465, B => n5470, Z => n5484);
   U5091 : AO2 port map( A => n5486, B => n5487, C => n5488, D => n5489, Z => 
                           n5481);
   U5092 : NR2 port map( A => n5490, B => n5491, Z => n5488);
   U5093 : NR2 port map( A => n5492, B => n5493, Z => n5486);
   U5094 : OR4 port map( A => n5494, B => n5495, C => n5496, D => n5497, Z => 
                           n5420);
   U5095 : AO4 port map( A => n5498, B => n5435, C => n5499, D => n5444, Z => 
                           n5497);
   U5096 : MUX21L port map( A => n5473, B => n5431, S => n4677, Z => n5496);
   U5097 : AO4 port map( A => n5500, B => n5479, C => n5501, D => n4643, Z => 
                           n5495);
   U5098 : AO4 port map( A => n5502, B => n5503, C => n5440, D => n5504, Z => 
                           n5494);
   U5099 : ND2 port map( A => n5505, B => n5506, Z => n5504);
   U5100 : ND2 port map( A => v_RAM_OUT0_13_port, B => n4398, Z => n5503);
   U5101 : AO7 port map( A => n5507, B => n5009, C => n5508, Z => n4183);
   U5102 : AO2 port map( A => n5418, B => n4620, C => n7813, D => n5419, Z => 
                           n5508);
   U5103 : AN2 port map( A => n5509, B => n5510, Z => n4620);
   U5104 : AO7 port map( A => n5511, B => n5512, C => n5513, Z => n5510);
   U5105 : AO3 port map( A => n5473, B => n5514, C => n5515, D => n5516, Z => 
                           n5512);
   U5106 : MUX21L port map( A => n5517, B => n5518, S => n5519, Z => n5516);
   U5107 : NR2 port map( A => n5442, B => n4649, Z => n5518);
   U5108 : NR2 port map( A => n5520, B => n5444, Z => n5517);
   U5109 : MUX21L port map( A => n5483, B => n5476, S => n5521, Z => n5515);
   U5110 : AO3 port map( A => n4357, B => n5505, C => n5522, D => n5523, Z => 
                           n5511);
   U5111 : AO2 port map( A => n5524, B => n5485, C => n5525, D => n5526, Z => 
                           n5523);
   U5112 : AO7 port map( A => n5527, B => n5528, C => n5477, Z => n5522);
   U5113 : MUX21L port map( A => n5529, B => n5530, S => n4361, Z => n5509);
   U5114 : AO4 port map( A => n5531, B => n4661, C => n5532, D => n5533, Z => 
                           n5530);
   U5115 : AO1 port map( A => n5534, B => n5461, C => n5535, D => n5536, Z => 
                           n5532);
   U5116 : AO6 port map( A => n5502, B => n5537, C => n5463, Z => n5536);
   U5117 : AO4 port map( A => n5436, B => n5456, C => n5432, D => n5538, Z => 
                           n5535);
   U5118 : ND2 port map( A => n5537, B => n5539, Z => n5534);
   U5119 : AO1 port map( A => n4678, B => n5540, C => n5541, D => n5542, Z => 
                           n5531);
   U5120 : NR2 port map( A => n5463, B => n5543, Z => n5542);
   U5121 : AO3 port map( A => n5464, B => n5505, C => n5544, D => n5545, Z => 
                           n5541);
   U5122 : AO7 port map( A => n5546, B => n5547, C => n5548, Z => n5544);
   U5123 : AO6 port map( A => n5549, B => n5550, C => n5551, Z => n5529);
   U5124 : AO4 port map( A => n5552, B => n4661, C => n5553, D => n5554, Z => 
                           n5551);
   U5125 : ND2 port map( A => n4665, B => n5545, Z => n5554);
   U5126 : ND2 port map( A => n5555, B => n5469, Z => n5545);
   U5127 : MUX21L port map( A => n5464, B => n5556, S => n5557, Z => n5553);
   U5128 : NR2 port map( A => n5548, B => n5558, Z => n5556);
   U5129 : AO6 port map( A => n5539, B => n4644, C => n5456, Z => n5558);
   U5130 : AO1 port map( A => n5559, B => n5548, C => n5560, D => n5561, Z => 
                           n5552);
   U5131 : AO4 port map( A => n5464, B => n5562, C => n5563, D => n5456, Z => 
                           n5560);
   U5132 : NR2 port map( A => n5564, B => n5459, Z => n5563);
   U5133 : NR2 port map( A => n5555, B => n5493, Z => n5559);
   U5134 : AO1 port map( A => n5565, B => n5525, C => n5566, D => n5567, Z => 
                           n5550);
   U5135 : AO4 port map( A => n5568, B => n5569, C => n5437, D => n5480, Z => 
                           n5567);
   U5136 : ND2 port map( A => n5521, B => n5465, Z => n5480);
   U5137 : ND2 port map( A => v_RAM_OUT0_13_port, B => n4357, Z => n5569);
   U5138 : IV port map( A => n5547, Z => n5568);
   U5139 : AO4 port map( A => n5473, B => n5446, C => n5502, D => n5435, Z => 
                           n5566);
   U5140 : IV port map( A => n5570, Z => n5565);
   U5141 : AO1 port map( A => n4676, B => n5485, C => n5571, D => n4397, Z => 
                           n5549);
   U5142 : AO4 port map( A => n5431, B => n5572, C => n5573, D => n5440, Z => 
                           n5571);
   U5143 : NR2 port map( A => n5574, B => n5498, Z => n5573);
   U5144 : AO7 port map( A => n5575, B => n5009, C => n5576, Z => n4182);
   U5145 : AO2 port map( A => n5418, B => n4624, C => n7883, D => n5419, Z => 
                           n5576);
   U5146 : AN2 port map( A => n5577, B => n5578, Z => n4624);
   U5147 : AO3 port map( A => n5579, B => n5580, C => n4353, D => n5513, Z => 
                           n5578);
   U5148 : IV port map( A => n5581, Z => n5580);
   U5149 : AO6 port map( A => n5461, B => n4645, C => n5582, Z => n5581);
   U5150 : AO4 port map( A => n5432, B => n5583, C => n5584, D => n5463, Z => 
                           n5579);
   U5151 : NR2 port map( A => n5490, B => n5460, Z => n5584);
   U5152 : MUX21L port map( A => n5585, B => n5586, S => n4361, Z => n5577);
   U5153 : AO3 port map( A => n5587, B => n5533, C => n5588, D => n5589, Z => 
                           n5586);
   U5154 : ND2 port map( A => n4667, B => n5590, Z => n5589);
   U5155 : AO3 port map( A => n5464, B => n5591, C => n5592, D => n5593, Z => 
                           n5590);
   U5156 : AO6 port map( A => n5540, B => n4674, C => n5561, Z => n5593);
   U5157 : MUX21L port map( A => n5469, B => n5594, S => n5595, Z => n5592);
   U5158 : NR2 port map( A => n5574, B => n5432, Z => n5594);
   U5159 : AO3 port map( A => n5463, B => n5572, C => n5596, D => n5597, Z => 
                           n5588);
   U5160 : AO6 port map( A => n4678, B => n5548, C => n4661, Z => n5597);
   U5161 : AO2 port map( A => n5501, B => n5461, C => n5540, D => n5598, Z => 
                           n5596);
   U5162 : ND2 port map( A => n5446, B => n5478, Z => n5598);
   U5163 : IV port map( A => n5599, Z => n5572);
   U5164 : AO1 port map( A => n4674, B => n5461, C => n5600, D => n5601, Z => 
                           n5587);
   U5165 : AO4 port map( A => n5432, B => n5602, C => n5603, D => n5456, Z => 
                           n5600);
   U5166 : AO3 port map( A => n5604, B => n4397, C => n5605, D => n5606, Z => 
                           n5585);
   U5167 : AO3 port map( A => n5464, B => n5607, C => n5453, D => n5608, Z => 
                           n5606);
   U5168 : AO6 port map( A => n4673, B => n5469, C => n5609, Z => n5608);
   U5169 : AO4 port map( A => n5456, B => n5610, C => n4357, D => n5611, Z => 
                           n5609);
   U5170 : ND2 port map( A => n4677, B => n5447, Z => n5607);
   U5171 : ND2 port map( A => n4665, B => n5612, Z => n5605);
   U5172 : AO3 port map( A => n4352, B => n4398, C => n5613, D => n5614, Z => 
                           n5612);
   U5173 : AO2 port map( A => n5520, B => n4357, C => n5469, D => n5611, Z => 
                           n5614);
   U5174 : MUX21H port map( A => n5434, B => n4674, S => n5548, Z => n5613);
   U5175 : NR4 port map( A => n5615, B => n5616, C => n5617, D => n5618, Z => 
                           n5604);
   U5176 : AO6 port map( A => n5431, B => n5473, C => n5521, Z => n5618);
   U5177 : EON1 port map( A => n5444, B => n5471, C => n5619, D => n5475, Z => 
                           n5616);
   U5178 : ND2 port map( A => n5620, B => n5621, Z => n5615);
   U5179 : EO1 port map( A => n5476, B => n4674, C => n5435, D => n5622, Z => 
                           n5621);
   U5180 : AO2 port map( A => n5524, B => n5485, C => n5525, D => n5623, Z => 
                           n5620);
   U5181 : AO7 port map( A => n5624, B => n5009, C => n5625, Z => n4181);
   U5182 : AO2 port map( A => n5418, B => n4627, C => n7812, D => n5419, Z => 
                           n5625);
   U5183 : MUX21L port map( A => n5626, B => n5627, S => n4361, Z => n4627);
   U5184 : AO1 port map( A => n4667, B => n5628, C => n5629, D => n5630, Z => 
                           n5627);
   U5185 : AO1 port map( A => n5520, B => n5461, C => n5631, D => n5632, Z => 
                           n5630);
   U5186 : AO4 port map( A => n5463, B => n5633, C => n5634, D => n5456, Z => 
                           n5632);
   U5187 : AO6 port map( A => v_RAM_OUT0_11_port, B => n4352, C => n5493, Z => 
                           n5634);
   U5188 : AO7 port map( A => n5432, B => n4674, C => n4665, Z => n5631);
   U5189 : AO4 port map( A => n5635, B => n4397, C => n5636, D => n4661, Z => 
                           n5629);
   U5190 : AO1 port map( A => n5548, B => n5538, C => n5637, D => n5638, Z => 
                           n5636);
   U5191 : AN3 port map( A => n5461, B => n5537, C => n5502, Z => n5638);
   U5192 : AO4 port map( A => n5456, B => n5543, C => n5463, D => n5468, Z => 
                           n5637);
   U5193 : IV port map( A => n5500, Z => n5468);
   U5194 : IV port map( A => n5493, Z => n5543);
   U5195 : NR4 port map( A => n5639, B => n5640, C => n5525, D => n5641, Z => 
                           n5635);
   U5196 : AN3 port map( A => n5539, B => n5611, C => n5485, Z => n5641);
   U5197 : AN3 port map( A => n5499, B => n4353, C => n4398, Z => n5640);
   U5198 : AO4 port map( A => n5464, B => n5470, C => n5622, D => n4649, Z => 
                           n5639);
   U5199 : AO3 port map( A => n5463, B => n5642, C => n5643, D => n5644, Z => 
                           n5628);
   U5200 : MUX21L port map( A => n5548, B => n5540, S => n5524, Z => n5644);
   U5201 : IV port map( A => n5561, Z => n5643);
   U5202 : AO1 port map( A => n5453, B => n5645, C => n5646, D => n5647, Z => 
                           n5626);
   U5203 : AN4 port map( A => n5648, B => n5649, C => n4665, D => n5650, Z => 
                           n5647);
   U5204 : AO2 port map( A => n5548, B => n5460, C => n5469, D => n5475, Z => 
                           n5650);
   U5205 : AO2 port map( A => n5461, B => n5546, C => n5570, D => n5540, Z => 
                           n5649);
   U5206 : ND2 port map( A => n5561, B => n5651, Z => n5648);
   U5207 : NR2 port map( A => n5470, B => n5463, Z => n5561);
   U5208 : AO4 port map( A => n5652, B => n5653, C => n5654, D => n4397, Z => 
                           n5646);
   U5209 : AO1 port map( A => n5655, B => n5656, C => n5657, D => n5658, Z => 
                           n5654);
   U5210 : NR3 port map( A => n5475, B => n5430, C => n5473, Z => n5658);
   U5211 : NR3 port map( A => n5659, B => n4645, C => n5479, Z => n5657);
   U5212 : ND2 port map( A => n5431, B => n5660, Z => n5655);
   U5213 : OR3 port map( A => n4398, B => v_RAM_OUT0_13_port, C => n5447, Z => 
                           n5660);
   U5214 : AO1 port map( A => n5469, B => n5661, C => n5662, D => n5663, Z => 
                           n5652);
   U5215 : AN3 port map( A => n5540, B => n5562, C => n5433, Z => n5663);
   U5216 : AO4 port map( A => n5432, B => n5664, C => n5464, D => n5665, Z => 
                           n5662);
   U5217 : ND2 port map( A => n5526, B => n5557, Z => n5665);
   U5218 : ND2 port map( A => n5539, B => n5611, Z => n5664);
   U5219 : ND2 port map( A => n5591, B => n5526, Z => n5661);
   U5220 : AO3 port map( A => n5464, B => n5666, C => n5667, D => n5668, Z => 
                           n5645);
   U5221 : AO2 port map( A => n5669, B => n5540, C => n5491, D => n5469, Z => 
                           n5668);
   U5222 : ND3 port map( A => n5447, B => n4677, C => n5548, Z => n5667);
   U5223 : IV port map( A => n5670, Z => n5447);
   U5224 : AO7 port map( A => n5671, B => n5009, C => n5672, Z => n4180);
   U5225 : AO2 port map( A => n5418, B => n4630, C => n7811, D => n5419, Z => 
                           n5672);
   U5226 : IV port map( A => n5673, Z => n4630);
   U5227 : AO3 port map( A => n5674, B => n5675, C => n5676, D => n5677, Z => 
                           n5673);
   U5228 : AO2 port map( A => n5421, B => n5678, C => v_RAM_OUT0_9_port, D => 
                           n5679, Z => n5677);
   U5229 : AO4 port map( A => n5680, B => n5533, C => n5681, D => n4661, Z => 
                           n5679);
   U5230 : AO6 port map( A => n5548, B => n5656, C => n5682, Z => n5681);
   U5231 : AO4 port map( A => n5456, B => n5462, C => n5683, D => n5684, Z => 
                           n5682);
   U5232 : IV port map( A => n4671, Z => n5684);
   U5233 : AO6 port map( A => n5685, B => n4357, C => n5461, Z => n5683);
   U5234 : AO1 port map( A => n5548, B => n5633, C => n5686, D => n5687, Z => 
                           n5680);
   U5235 : AO6 port map( A => n5595, B => n5433, C => n5464, Z => n5687);
   U5236 : IV port map( A => n4645, Z => n5595);
   U5237 : AO4 port map( A => n5441, B => n5463, C => n5456, D => n5539, Z => 
                           n5686);
   U5238 : IV port map( A => n5455, Z => n5633);
   U5239 : ND4 port map( A => n5688, B => n5689, C => n5690, D => n5691, Z => 
                           n5678);
   U5240 : AO2 port map( A => n5476, B => n5692, C => n5483, D => n5693, Z => 
                           n5691);
   U5241 : ND2 port map( A => n5623, B => n5656, Z => n5693);
   U5242 : ND2 port map( A => n5465, B => n5583, Z => n5692);
   U5243 : IV port map( A => n5546, Z => n5583);
   U5244 : AO2 port map( A => n5669, B => n5477, C => n5489, D => n5514, Z => 
                           n5690);
   U5245 : MUX21L port map( A => n5485, B => n5694, S => n5611, Z => n5689);
   U5246 : NR2 port map( A => n5695, B => n5444, Z => n5694);
   U5247 : AO2 port map( A => n4646, B => n5436, C => n4676, D => n5525, Z => 
                           n5688);
   U5248 : ND4 port map( A => n5696, B => n5697, C => n5698, D => n5699, Z => 
                           n5676);
   U5249 : AO1 port map( A => n5500, B => n5483, C => n5700, D => n4647, Z => 
                           n5699);
   U5250 : IV port map( A => n5513, Z => n4647);
   U5251 : AO4 port map( A => n5701, B => n5437, C => n5702, D => n5444, Z => 
                           n5700);
   U5252 : AN2 port map( A => n5478, B => n4677, Z => n5702);
   U5253 : NR2 port map( A => n5519, B => n5493, Z => n5500);
   U5254 : AO1 port map( A => n5703, B => n5525, C => n5704, D => n5617, Z => 
                           n5698);
   U5255 : NR2 port map( A => n5465, B => n5473, Z => n5617);
   U5256 : NR2 port map( A => v_RAM_OUT0_11_port, B => n5520, Z => n5703);
   U5257 : ND3 port map( A => n5591, B => n5526, C => n5485, Z => n5697);
   U5258 : OR3 port map( A => n5695, B => n5441, C => n5435, Z => n5696);
   U5259 : AO3 port map( A => n5599, B => n5431, C => n5705, D => n4639, Z => 
                           n5675);
   U5260 : AO7 port map( A => v_RAM_OUT0_8_port, B => n4408, C => n5485, Z => 
                           n5705);
   U5261 : NR2 port map( A => n5547, B => n5528, Z => n5599);
   U5262 : AO3 port map( A => n5446, B => n5706, C => n5707, D => n5708, Z => 
                           n5674);
   U5263 : AO2 port map( A => n5498, B => n4646, C => n5525, D => n5709, Z => 
                           n5708);
   U5264 : ND2 port map( A => n5433, B => n5537, Z => n5709);
   U5265 : AO3 port map( A => n5463, B => n5602, C => n5710, D => n5711, Z => 
                           n5707);
   U5266 : AO6 port map( A => n5701, B => n5540, C => n4353, Z => n5711);
   U5267 : AO2 port map( A => n5712, B => n5656, C => n5548, D => n5685, Z => 
                           n5710);
   U5268 : ND2 port map( A => n5478, B => n5539, Z => n5685);
   U5269 : NR2 port map( A => n5499, B => n5464, Z => n5712);
   U5270 : IV port map( A => n5490, Z => n5446);
   U5271 : AO7 port map( A => n5713, B => n5009, C => n5714, Z => n4179);
   U5272 : AO2 port map( A => n5418, B => n4769, C => n7810, D => n5419, Z => 
                           n5714);
   U5273 : AO1 port map( A => n4634, B => v_RAM_OUT0_9_port, C => n5715, D => 
                           n5716, Z => n4769);
   U5274 : AO1 port map( A => v_RAM_OUT0_13_port, B => n5717, C => n5718, D => 
                           n5719, Z => n5716);
   U5275 : AO7 port map( A => n4649, B => n4651, C => n5513, Z => n5719);
   U5276 : MUX21L port map( A => n5720, B => v_RAM_OUT0_12_port, S => n5519, Z 
                           => n4651);
   U5277 : NR2 port map( A => v_RAM_OUT0_12_port, B => n5520, Z => n5720);
   U5278 : ND2 port map( A => n4353, B => n4357, Z => n4649);
   U5279 : AO4 port map( A => n5473, B => n5721, C => n5462, D => n4643, Z => 
                           n5718);
   U5280 : IV port map( A => n5485, Z => n4643);
   U5281 : ND2 port map( A => n4644, B => n5521, Z => n5462);
   U5282 : IV port map( A => n5491, Z => n4644);
   U5283 : NR2 port map( A => n5695, B => n5722, Z => n5721);
   U5284 : IV port map( A => n4640, Z => n5717);
   U5285 : AO3 port map( A => n5464, B => n5723, C => n5724, D => n5725, Z => 
                           n4640);
   U5286 : ND3 port map( A => n5591, B => n5526, C => n5540, Z => n5725);
   U5287 : ND2 port map( A => n5726, B => n5465, Z => n5724);
   U5288 : AO7 port map( A => n5430, B => n5463, C => n5432, Z => n5726);
   U5289 : NR2 port map( A => n5727, B => n4638, Z => n5715);
   U5290 : AN4 port map( A => n5728, B => n5729, C => n5730, D => n5731, Z => 
                           n4638);
   U5291 : AO1 port map( A => n4646, B => n5732, C => n5733, D => n5734, Z => 
                           n5731);
   U5292 : AO6 port map( A => n5431, B => n5435, C => n5433, Z => n5734);
   U5293 : AO6 port map( A => n5440, B => n5437, C => n5610, Z => n5733);
   U5294 : ND2 port map( A => n5478, B => n5526, Z => n5732);
   U5295 : IV port map( A => n5735, Z => n5526);
   U5296 : AO2 port map( A => n5525, B => n5736, C => n5547, D => n5619, Z => 
                           n5730);
   U5297 : ND2 port map( A => n5440, B => n5444, Z => n5619);
   U5298 : ND2 port map( A => n5465, B => n5656, Z => n5736);
   U5299 : AO2 port map( A => n5527, B => n5477, C => n5528, D => n5487, Z => 
                           n5729);
   U5300 : AO2 port map( A => n5476, B => v_RAM_OUT0_11_port, C => n5460, D => 
                           n5485, Z => n5728);
   U5301 : IV port map( A => n4639, Z => n5727);
   U5302 : AO3 port map( A => n5737, B => n5533, C => n5738, D => n5739, Z => 
                           n4634);
   U5303 : ND3 port map( A => n5740, B => n5453, C => n5741, Z => n5739);
   U5304 : AO1 port map( A => n5548, B => n5742, C => n5651, D => n5743, Z => 
                           n5741);
   U5305 : AO6 port map( A => n5465, B => n5506, C => n5456, Z => n5743);
   U5306 : ND2 port map( A => n5434, B => n5610, Z => n5742);
   U5307 : AO2 port map( A => n5603, B => n5469, C => n5564, D => n4398, Z => 
                           n5740);
   U5308 : IV port map( A => n5744, Z => n5603);
   U5309 : ND4 port map( A => n5745, B => n5746, C => n5747, D => n5748, Z => 
                           n5738);
   U5310 : AO1 port map( A => n5525, B => n5499, C => n5749, D => n4397, Z => 
                           n5748);
   U5311 : AO4 port map( A => n5695, B => n5473, C => n5440, D => n5514, Z => 
                           n5749);
   U5312 : AO2 port map( A => n5485, B => n5505, C => n5442, D => n5477, Z => 
                           n5747);
   U5313 : IV port map( A => n5527, Z => n5505);
   U5314 : NR2 port map( A => n5623, B => v_RAM_OUT0_8_port, Z => n5527);
   U5315 : AO7 port map( A => n5476, B => n5489, C => n5750, Z => n5746);
   U5316 : AO2 port map( A => n5751, B => n5487, C => n5752, D => n5564, Z => 
                           n5745);
   U5317 : NR2 port map( A => v_RAM_OUT0_13_port, B => n4398, Z => n5752);
   U5318 : AN2 port map( A => n5537, B => n5539, Z => n5751);
   U5319 : AO1 port map( A => n5753, B => n5548, C => n5754, D => n5651, Z => 
                           n5737);
   U5320 : NR2 port map( A => n5478, B => n5464, Z => n5651);
   U5321 : AO4 port map( A => n5456, B => n5519, C => n5755, D => n5463, Z => 
                           n5754);
   U5322 : NR2 port map( A => n5750, B => n5574, Z => n5755);
   U5323 : NR2 port map( A => n5670, B => n5490, Z => n5753);
   U5324 : AO7 port map( A => n5756, B => n5009, C => n5757, Z => n4178);
   U5325 : AO2 port map( A => n5418, B => n4654, C => n7809, D => n5419, Z => 
                           n5757);
   U5326 : IV port map( A => n5758, Z => n4654);
   U5327 : AO3 port map( A => n5759, B => n5760, C => n5761, D => n5762, Z => 
                           n5758);
   U5328 : AO2 port map( A => n5421, B => n5763, C => v_RAM_OUT0_9_port, D => 
                           n5764, Z => n5762);
   U5329 : AO3 port map( A => n5765, B => n4661, C => n5766, D => n5767, Z => 
                           n5764);
   U5330 : OR3 port map( A => n5472, B => n5432, C => n5471, Z => n5767);
   U5331 : NR2 port map( A => n5453, B => n4665, Z => n5472);
   U5332 : AO7 port map( A => n5582, B => n5768, C => n4665, Z => n5766);
   U5333 : AO4 port map( A => n5464, B => n5434, C => n5501, D => n5463, Z => 
                           n5768);
   U5334 : NR2 port map( A => n5441, B => n5735, Z => n5501);
   U5335 : AO3 port map( A => n5432, B => n5465, C => n5769, D => n5770, Z => 
                           n5582);
   U5336 : ND3 port map( A => n5611, B => n5656, C => n5540, Z => n5770);
   U5337 : ND2 port map( A => n5493, B => n5461, Z => n5769);
   U5338 : IV port map( A => n5441, Z => n5465);
   U5339 : IV port map( A => n5453, Z => n4661);
   U5340 : AO1 port map( A => n5723, B => n5540, C => n5771, D => n5772, Z => 
                           n5765);
   U5341 : AO6 port map( A => n5591, B => n5506, C => n5463, Z => n5772);
   U5342 : IV port map( A => n5528, Z => n5506);
   U5343 : AO4 port map( A => n5432, B => n5562, C => n5455, D => n5464, Z => 
                           n5771);
   U5344 : AO3 port map( A => n5622, B => n5431, C => n5773, D => n5774, Z => 
                           n5763);
   U5345 : AO1 port map( A => n5775, B => n5557, C => n5776, D => n5777, Z => 
                           n5774);
   U5346 : AO6 port map( A => n5436, B => n5610, C => n5440, Z => n5777);
   U5347 : IV port map( A => n5483, Z => n5440);
   U5348 : AO4 port map( A => n5444, B => n5602, C => n5438, D => n5473, Z => 
                           n5776);
   U5349 : NR2 port map( A => n5490, B => n5722, Z => n5438);
   U5350 : IV port map( A => n5475, Z => n5602);
   U5351 : IV port map( A => n5487, Z => n5444);
   U5352 : AO7 port map( A => n5735, B => n5479, C => n5437, Z => n5775);
   U5353 : AO2 port map( A => n5493, B => n5477, C => n4676, D => n5485, Z => 
                           n5773);
   U5354 : NR2 port map( A => n5735, B => n5460, Z => n5622);
   U5355 : NR2 port map( A => n5519, B => n4352, Z => n5735);
   U5356 : NR2 port map( A => n4361, B => n4397, Z => n5421);
   U5357 : AO3 port map( A => n5431, B => n5478, C => n5513, D => n5778, Z => 
                           n5761);
   U5358 : AO1 port map( A => n4676, B => n5779, C => n5780, D => n5781, Z => 
                           n5778);
   U5359 : NR3 port map( A => n5574, B => n5498, C => n5479, Z => n5781);
   U5360 : AO1 port map( A => n5540, B => v_RAM_OUT0_11_port, C => n5782, D => 
                           n4353, Z => n5780);
   U5361 : AO3 port map( A => n5464, B => n5744, C => n5783, D => n5784, Z => 
                           n5782);
   U5362 : ND3 port map( A => n5519, B => n5656, C => n5469, Z => n5784);
   U5363 : IV port map( A => n5695, Z => n5656);
   U5364 : AO7 port map( A => n5659, B => n5460, C => n5548, Z => n5783);
   U5365 : AO7 port map( A => n5591, B => n5706, C => n5473, Z => n5779);
   U5366 : NR2 port map( A => n4397, B => v_RAM_OUT0_9_port, Z => n5513);
   U5367 : AO3 port map( A => n5479, B => n5642, C => n4639, D => n5785, Z => 
                           n5760);
   U5368 : AO2 port map( A => n5483, B => n5666, C => n5485, D => n4674, Z => 
                           n5785);
   U5369 : NR2 port map( A => n5456, B => v_RAM_OUT0_13_port, Z => n5485);
   U5370 : NR2 port map( A => n4353, B => n5456, Z => n5483);
   U5371 : NR2 port map( A => v_RAM_OUT0_9_port, B => v_RAM_OUT0_15_port, Z => 
                           n4639);
   U5372 : ND4 port map( A => n5786, B => n5787, C => n5788, D => n5789, Z => 
                           n5759);
   U5373 : AO2 port map( A => n5487, B => n5570, C => n5455, D => n4646, Z => 
                           n5789);
   U5374 : NR2 port map( A => n5546, B => n5670, Z => n5455);
   U5375 : NR2 port map( A => n5492, B => v_RAM_OUT0_8_port, Z => n5670);
   U5376 : ND2 port map( A => n5557, B => n5610, Z => n5570);
   U5377 : IV port map( A => n5520, Z => n5610);
   U5378 : NR2 port map( A => n4352, B => n5492, Z => n5520);
   U5379 : NR2 port map( A => n5463, B => n4353, Z => n5487);
   U5380 : OR3 port map( A => n5441, B => n5442, C => n5435, Z => n5788);
   U5381 : IV port map( A => n5477, Z => n5435);
   U5382 : NR2 port map( A => n4353, B => n5464, Z => n5477);
   U5383 : IV port map( A => n5704, Z => n5787);
   U5384 : NR3 port map( A => n5750, B => n5546, C => n5431, Z => n5704);
   U5385 : OR3 port map( A => n5491, B => n5490, C => n5437, Z => n5786);
   U5386 : IV port map( A => n5476, Z => n5437);
   U5387 : NR2 port map( A => n5432, B => n4353, Z => n5476);
   U5388 : AO7 port map( A => n5790, B => n5009, C => n5791, Z => n4177);
   U5389 : AO2 port map( A => n5418, B => n4774, C => n7808, D => n5419, Z => 
                           n5791);
   U5390 : MUX21L port map( A => n5792, B => n4660, S => n4361, Z => n4774);
   U5391 : AO3 port map( A => n5793, B => n5533, C => n5794, D => n5795, Z => 
                           n4660);
   U5392 : AO2 port map( A => v_RAM_OUT0_15_port, B => n5796, C => n4667, D => 
                           n5797, Z => n5795);
   U5393 : AO3 port map( A => n5456, B => n5538, C => n5798, D => n5799, Z => 
                           n5797);
   U5394 : AO2 port map( A => n5469, B => n5514, C => n5548, D => n5436, Z => 
                           n5799);
   U5395 : ND2 port map( A => n5478, B => n5471, Z => n5514);
   U5396 : AO7 port map( A => n5490, B => n5491, C => n5461, Z => n5798);
   U5397 : AO7 port map( A => n5524, B => n5479, C => n5800, Z => n5796);
   U5398 : EO1 port map( A => n5801, B => n5802, C => n5538, D => n5431, Z => 
                           n5800);
   U5399 : ND2 port map( A => n5434, B => n4677, Z => n5538);
   U5400 : IV port map( A => n5442, Z => n4677);
   U5401 : AO7 port map( A => n5537, B => n5706, C => n5473, Z => n5801);
   U5402 : IV port map( A => n4646, Z => n5473);
   U5403 : ND2 port map( A => v_RAM_OUT0_10_port, B => n4353, Z => n5706);
   U5404 : IV port map( A => n5459, Z => n5537);
   U5405 : IV port map( A => n5525, Z => n5479);
   U5406 : NR2 port map( A => n5464, B => v_RAM_OUT0_13_port, Z => n5525);
   U5407 : NR2 port map( A => n5803, B => n5460, Z => n5524);
   U5408 : NR2 port map( A => n5611, B => v_RAM_OUT0_8_port, Z => n5460);
   U5409 : AO3 port map( A => n5441, B => n5456, C => n5453, D => n5804, Z => 
                           n5794);
   U5410 : AO1 port map( A => n5805, B => n5461, C => n4642, D => n5601, Z => 
                           n5804);
   U5411 : AN3 port map( A => n5433, B => n5642, C => n5469, Z => n5601);
   U5412 : IV port map( A => n5750, Z => n5642);
   U5413 : NR2 port map( A => v_RAM_OUT0_8_port, B => n5701, Z => n5750);
   U5414 : IV port map( A => n5574, Z => n5433);
   U5415 : NR2 port map( A => n4352, B => v_RAM_OUT0_11_port, Z => n5574);
   U5416 : NR2 port map( A => n5521, B => n4357, Z => n4642);
   U5417 : IV port map( A => n5564, Z => n5521);
   U5418 : NR2 port map( A => n5434, B => n4352, Z => n5564);
   U5419 : ND2 port map( A => n5471, B => n5562, Z => n5805);
   U5420 : IV port map( A => n5498, Z => n5562);
   U5421 : NR2 port map( A => n5434, B => v_RAM_OUT0_8_port, Z => n5498);
   U5422 : IV port map( A => n5701, Z => n5434);
   U5423 : IV port map( A => n5430, Z => n5471);
   U5424 : NR2 port map( A => v_RAM_OUT0_8_port, B => v_RAM_OUT0_11_port, Z => 
                           n5441);
   U5425 : AO1 port map( A => n5469, B => n5539, C => n5806, D => n5807, Z => 
                           n5793);
   U5426 : NR2 port map( A => n5464, B => n5669, Z => n5807);
   U5427 : AO4 port map( A => v_RAM_OUT0_11_port, B => n5432, C => n5557, D => 
                           n5456, Z => n5806);
   U5428 : NR2 port map( A => n5808, B => n5809, Z => n5792);
   U5429 : AO4 port map( A => n5653, B => n4668, C => n5533, D => n4666, Z => 
                           n5809);
   U5430 : AO3 port map( A => n5723, B => n5432, C => n5810, D => n5811, Z => 
                           n4666);
   U5431 : EO1 port map( A => n5546, B => n5540, C => n5669, D => n5464, Z => 
                           n5811);
   U5432 : NR2 port map( A => n5442, B => n5547, Z => n5669);
   U5433 : NR2 port map( A => v_RAM_OUT0_8_port, B => n5499, Z => n5547);
   U5434 : NR2 port map( A => n4366, B => n4352, Z => n5546);
   U5435 : AO7 port map( A => n5695, B => n5491, C => n5469, Z => n5810);
   U5436 : NR2 port map( A => n5491, B => n5493, Z => n5723);
   U5437 : NR2 port map( A => n4352, B => n5499, Z => n5493);
   U5438 : IV port map( A => n4665, Z => n5533);
   U5439 : NR2 port map( A => v_RAM_OUT0_15_port, B => v_RAM_OUT0_13_port, Z =>
                           n4665);
   U5440 : AO3 port map( A => n5812, B => n5456, C => n5813, D => n5814, Z => 
                           n4668);
   U5441 : AO2 port map( A => n5744, B => n5461, C => n5469, D => n5539, Z => 
                           n5814);
   U5442 : ND2 port map( A => v_RAM_OUT0_8_port, B => n5519, Z => n5539);
   U5443 : ND2 port map( A => n5502, B => n5478, Z => n5744);
   U5444 : ND2 port map( A => n4352, B => n4366, Z => n5478);
   U5445 : IV port map( A => n5803, Z => n5502);
   U5446 : AO7 port map( A => n5490, B => n5459, C => v_RAM_OUT0_10_port, Z => 
                           n5813);
   U5447 : NR2 port map( A => n5557, B => v_RAM_OUT0_8_port, Z => n5459);
   U5448 : NR2 port map( A => n5623, B => n4352, Z => n5490);
   U5449 : IV port map( A => n5492, Z => n5623);
   U5450 : NR2 port map( A => n5695, B => n5475, Z => n5812);
   U5451 : NR2 port map( A => v_RAM_OUT0_8_port, B => n5555, Z => n5475);
   U5452 : NR2 port map( A => n4352, B => n5701, Z => n5695);
   U5453 : IV port map( A => n4667, Z => n5653);
   U5454 : NR2 port map( A => n4353, B => n4397, Z => n4667);
   U5455 : EON1 port map( A => n5815, B => n4397, C => n5816, D => n5453, Z => 
                           n5808);
   U5456 : NR2 port map( A => n4353, B => v_RAM_OUT0_15_port, Z => n5453);
   U5457 : AO7 port map( A => n5432, B => n5442, C => n5817, Z => n5816);
   U5458 : AO2 port map( A => n5802, B => n4672, C => n5469, D => n4678, Z => 
                           n5817);
   U5459 : NR2 port map( A => n5430, B => n4645, Z => n4678);
   U5460 : NR2 port map( A => n5611, B => n4352, Z => n5430);
   U5461 : IV port map( A => n5555, Z => n5611);
   U5462 : IV port map( A => n4676, Z => n5802);
   U5463 : NR2 port map( A => n5803, B => n4645, Z => n4676);
   U5464 : NR2 port map( A => n5519, B => v_RAM_OUT0_8_port, Z => n4645);
   U5465 : IV port map( A => n5436, Z => n5519);
   U5466 : NR2 port map( A => n4352, B => n4408, Z => n5803);
   U5467 : AO1 port map( A => n4646, B => n5666, C => n5818, D => n5819, Z => 
                           n5815);
   U5468 : AN3 port map( A => n4672, B => n4353, C => n4671, Z => n5819);
   U5469 : NR2 port map( A => n5491, B => n5528, Z => n4671);
   U5470 : NR2 port map( A => n4352, B => n5557, Z => n5528);
   U5471 : IV port map( A => n5499, Z => n5557);
   U5472 : NR2 port map( A => n4408, B => v_RAM_OUT0_14_port, Z => n5499);
   U5473 : NR2 port map( A => n4366, B => v_RAM_OUT0_8_port, Z => n5491);
   U5474 : ND2 port map( A => n5464, B => n5456, Z => n4672);
   U5475 : IV port map( A => n5540, Z => n5456);
   U5476 : NR2 port map( A => n4398, B => n4357, Z => n5540);
   U5477 : IV port map( A => n5461, Z => n5464);
   U5478 : NR2 port map( A => v_RAM_OUT0_12_port, B => v_RAM_OUT0_10_port, Z =>
                           n5461);
   U5479 : NR2 port map( A => n5431, B => n4674, Z => n5818);
   U5480 : ND2 port map( A => n5470, B => n5591, Z => n4674);
   U5481 : IV port map( A => n5722, Z => n5591);
   U5482 : NR2 port map( A => v_RAM_OUT0_8_port, B => n5436, Z => n5722);
   U5483 : NR2 port map( A => n5555, B => n5701, Z => n5436);
   U5484 : NR2 port map( A => n4366, B => n4408, Z => n5701);
   U5485 : IV port map( A => n5659, Z => n5470);
   U5486 : NR2 port map( A => n4352, B => v_RAM_OUT0_14_port, Z => n5659);
   U5487 : IV port map( A => n5489, Z => n5431);
   U5488 : NR2 port map( A => n5463, B => v_RAM_OUT0_13_port, Z => n5489);
   U5489 : IV port map( A => n5469, Z => n5463);
   U5490 : NR2 port map( A => n4398, B => v_RAM_OUT0_10_port, Z => n5469);
   U5491 : IV port map( A => n4673, Z => n5666);
   U5492 : NR2 port map( A => n5442, B => n5492, Z => n4673);
   U5493 : NR2 port map( A => n4366, B => v_RAM_OUT0_11_port, Z => n5492);
   U5494 : NR2 port map( A => n4352, B => n5555, Z => n5442);
   U5495 : NR2 port map( A => v_RAM_OUT0_14_port, B => v_RAM_OUT0_11_port, Z =>
                           n5555);
   U5496 : NR2 port map( A => n5432, B => v_RAM_OUT0_13_port, Z => n4646);
   U5497 : IV port map( A => n5548, Z => n5432);
   U5498 : NR2 port map( A => n4357, B => v_RAM_OUT0_12_port, Z => n5548);
   U5499 : NR2 port map( A => n5384, B => n5419, Z => n5418);
   U5500 : NR2 port map( A => n5384, B => n4706, Z => n5419);
   U5501 : NR2 port map( A => n5385, B => n4526, Z => n4706);
   U5502 : OR3 port map( A => v_CALCULATION_CNTR_3_port, B => 
                           v_CALCULATION_CNTR_1_port, C => n4565, Z => n5385);
   U5503 : IV port map( A => n5820, Z => n5790);
   U5504 : AO7 port map( A => n5821, B => n5009, C => n5822, Z => n4176);
   U5505 : AO2 port map( A => n5823, B => n4681, C => n7875, D => n5824, Z => 
                           n5822);
   U5506 : IV port map( A => n5825, Z => n4681);
   U5507 : AO7 port map( A => n5826, B => n5827, C => n5828, Z => n5825);
   U5508 : MUX21L port map( A => n5829, B => n5830, S => n4395, Z => n5828);
   U5509 : AO3 port map( A => n5831, B => n5832, C => n5833, D => n5834, Z => 
                           n5830);
   U5510 : AO1 port map( A => n5835, B => n5836, C => n5837, D => n5838, Z => 
                           n5834);
   U5511 : AO6 port map( A => n5839, B => n5840, C => n5841, Z => n5838);
   U5512 : ND3 port map( A => v_RAM_OUT0_18_port, B => n5842, C => n5831, Z => 
                           n5840);
   U5513 : AN3 port map( A => n5843, B => n4358, C => n5844, Z => n5837);
   U5514 : EO1 port map( A => n5845, B => n5846, C => n4797, D => n5847, Z => 
                           n5833);
   U5515 : NR4 port map( A => n5848, B => n5849, C => n5850, D => n5851, Z => 
                           n5829);
   U5516 : AO4 port map( A => n5852, B => n5853, C => n4797, D => n5854, Z => 
                           n5851);
   U5517 : ND2 port map( A => n5855, B => n5856, Z => n5854);
   U5518 : ND2 port map( A => n5857, B => n4806, Z => n5853);
   U5519 : NR3 port map( A => n5858, B => v_RAM_OUT0_20_port, C => n5859, Z => 
                           n5850);
   U5520 : AO4 port map( A => n5860, B => n4805, C => n5861, D => n5862, Z => 
                           n5849);
   U5521 : AO1 port map( A => n5863, B => n5844, C => n5864, D => n5865, Z => 
                           n5860);
   U5522 : AO6 port map( A => n5866, B => n5867, C => n5858, Z => n5865);
   U5523 : AO4 port map( A => n5841, B => n4800, C => n5847, D => n5852, Z => 
                           n5864);
   U5524 : NR2 port map( A => n5868, B => n5869, Z => n5847);
   U5525 : AO3 port map( A => n5870, B => n5839, C => n5871, D => n5872, Z => 
                           n5848);
   U5526 : AO2 port map( A => n5873, B => n5874, C => n4801, D => n5875, Z => 
                           n5872);
   U5527 : AO3 port map( A => n4800, B => n5876, C => n5877, D => n5878, Z => 
                           n5875);
   U5528 : ND2 port map( A => n4820, B => n5879, Z => n5878);
   U5529 : OR3 port map( A => n5880, B => n5881, C => n5852, Z => n5877);
   U5530 : AO4 port map( A => n5882, B => n5858, C => n5852, D => n5883, Z => 
                           n5874);
   U5531 : MUX21L port map( A => n5884, B => n5846, S => n5885, Z => n5871);
   U5532 : NR4 port map( A => n5886, B => n5887, C => n5888, D => n5889, Z => 
                           n5826);
   U5533 : AO4 port map( A => n5890, B => n5856, C => n5891, D => n5892, Z => 
                           n5889);
   U5534 : AO4 port map( A => n5893, B => n5894, C => n5895, D => n5896, Z => 
                           n5888);
   U5535 : AO4 port map( A => n5897, B => n5898, C => n4358, D => n5899, Z => 
                           n5887);
   U5536 : MUX21L port map( A => n4822, B => n5900, S => n4363, Z => n5899);
   U5537 : AO4 port map( A => n5901, B => n5902, C => n5903, D => n5904, Z => 
                           n5886);
   U5538 : ND2 port map( A => n5905, B => n5906, Z => n5904);
   U5539 : AO7 port map( A => n5907, B => n5009, C => n5908, Z => n4175);
   U5540 : AO2 port map( A => n5823, B => n4686, C => n7889, D => n5824, Z => 
                           n5908);
   U5541 : MUX21L port map( A => n5909, B => n5910, S => n4395, Z => n4686);
   U5542 : AO1 port map( A => n5911, B => n5912, C => n5913, D => n5914, Z => 
                           n5910);
   U5543 : AO1 port map( A => n5857, B => n5915, C => n5916, D => n5917, Z => 
                           n5914);
   U5544 : AO4 port map( A => n5918, B => n5919, C => n5920, D => n5921, Z => 
                           n5917);
   U5545 : NR2 port map( A => n5882, B => n5900, Z => n5920);
   U5546 : AO7 port map( A => n5922, B => n4805, C => n5842, Z => n5916);
   U5547 : AO4 port map( A => n5923, B => n5858, C => n5924, D => n5852, Z => 
                           n5913);
   U5548 : AO1 port map( A => n5925, B => n4823, C => n5926, D => n5927, Z => 
                           n5924);
   U5549 : NR2 port map( A => v_RAM_OUT0_20_port, B => n5836, Z => n5927);
   U5550 : AO3 port map( A => n5928, B => n5929, C => n5930, D => n5931, Z => 
                           n5926);
   U5551 : ND3 port map( A => n5932, B => n5933, C => n4801, Z => n5930);
   U5552 : AO1 port map( A => n5934, B => n5873, C => n5935, D => n5936, Z => 
                           n5923);
   U5553 : AO4 port map( A => n5929, B => n5859, C => n5937, D => n4805, Z => 
                           n5935);
   U5554 : NR2 port map( A => n5938, B => n5900, Z => n5937);
   U5555 : NR2 port map( A => n5939, B => n5881, Z => n5934);
   U5556 : AO1 port map( A => n5939, B => n4801, C => n5940, D => n5941, Z => 
                           n5912);
   U5557 : NR2 port map( A => n4805, B => n5942, Z => n5941);
   U5558 : NR2 port map( A => n4808, B => n5943, Z => n5911);
   U5559 : MUX21L port map( A => n5929, B => n5918, S => n5944, Z => n5943);
   U5560 : MUX21L port map( A => n5945, B => n5946, S => n4403, Z => n5909);
   U5561 : AN3 port map( A => n5947, B => n5948, C => n5949, Z => n5946);
   U5562 : AO1 port map( A => n5950, B => n5951, C => n5952, D => n5953, Z => 
                           n5949);
   U5563 : NR4 port map( A => v_RAM_OUT0_18_port, B => v_RAM_OUT0_17_port, C =>
                           n5922, D => n4822, Z => n5953);
   U5564 : AO4 port map( A => n5903, B => n5954, C => n5896, D => n5955, Z => 
                           n5952);
   U5565 : NR2 port map( A => n5879, B => n5956, Z => n5950);
   U5566 : AO2 port map( A => n5957, B => n5958, C => n5959, D => n5960, Z => 
                           n5948);
   U5567 : EO1 port map( A => n5961, B => n5870, C => n5962, D => n5963, Z => 
                           n5947);
   U5568 : NR4 port map( A => n5964, B => n5965, C => n5966, D => n5967, Z => 
                           n5945);
   U5569 : AO4 port map( A => n5901, B => n4798, C => v_RAM_OUT0_17_port, D => 
                           n5866, Z => n5967);
   U5570 : MUX21L port map( A => n5896, B => n5968, S => n5855, Z => n5966);
   U5571 : AO6 port map( A => n5960, B => n5856, C => n5969, Z => n5968);
   U5572 : AO4 port map( A => n5867, B => n5898, C => n5970, D => n5971, Z => 
                           n5965);
   U5573 : AO6 port map( A => n5972, B => n5973, C => n5951, Z => n5971);
   U5574 : AO6 port map( A => n5974, B => n5859, C => n5890, Z => n5964);
   U5575 : AO7 port map( A => n5975, B => n5009, C => n5976, Z => n4174);
   U5576 : AO2 port map( A => n5823, B => n4689, C => n7890, D => n5824, Z => 
                           n5976);
   U5577 : MUX21H port map( A => n5977, B => n5978, S => v_RAM_OUT0_23_port, Z 
                           => n4689);
   U5578 : AO1 port map( A => n5979, B => n5980, C => n5981, D => n5982, Z => 
                           n5978);
   U5579 : AO4 port map( A => n5856, B => n5983, C => n5984, D => n5852, Z => 
                           n5982);
   U5580 : AO1 port map( A => n5891, B => n4801, C => n5985, D => n5986, Z => 
                           n5984);
   U5581 : AO7 port map( A => n5918, B => n5987, C => n5988, Z => n5986);
   U5582 : IV port map( A => n5936, Z => n5988);
   U5583 : AO4 port map( A => n5929, B => n5989, C => n5990, D => n4805, Z => 
                           n5985);
   U5584 : AO3 port map( A => n5991, B => n5858, C => n5992, D => n5993, Z => 
                           n5981);
   U5585 : AO2 port map( A => n5994, B => n5995, C => n5996, D => n5844, Z => 
                           n5993);
   U5586 : AO7 port map( A => n5846, B => n5884, C => n5938, Z => n5992);
   U5587 : AO1 port map( A => n5873, B => n4832, C => n5997, D => n5998, Z => 
                           n5991);
   U5588 : IV port map( A => n5999, Z => n5998);
   U5589 : AO6 port map( A => n6000, B => n5857, C => n6001, Z => n5999);
   U5590 : AO4 port map( A => n5921, B => n6002, C => n4805, D => n5883, Z => 
                           n5997);
   U5591 : AO1 port map( A => n5873, B => n6003, C => n6001, D => n6004, Z => 
                           n5980);
   U5592 : AO6 port map( A => n5932, B => n4804, C => n4805, Z => n6004);
   U5593 : ND2 port map( A => n5836, B => n6005, Z => n6003);
   U5594 : AO1 port map( A => n5857, B => n6006, C => n4800, D => n6007, Z => 
                           n5979);
   U5595 : NR2 port map( A => n5921, B => n6008, Z => n6007);
   U5596 : AO7 port map( A => n6009, B => n5858, C => n6010, Z => n5977);
   U5597 : MUX21L port map( A => n6011, B => n6012, S => n4403, Z => n6010);
   U5598 : NR4 port map( A => n6013, B => n6014, C => n6015, D => n6016, Z => 
                           n6012);
   U5599 : AO4 port map( A => n5893, B => n5890, C => n5883, D => n5963, Z => 
                           n6016);
   U5600 : MUX21L port map( A => n5892, B => n5898, S => n4832, Z => n6015);
   U5601 : AO4 port map( A => n5901, B => n6017, C => n6018, D => n5903, Z => 
                           n6014);
   U5602 : ND2 port map( A => n6019, B => n5974, Z => n6017);
   U5603 : EON1 port map( A => n6020, B => n5896, C => n6021, D => n5972, Z => 
                           n6013);
   U5604 : AO4 port map( A => n6022, B => n6023, C => n5890, D => n6008, Z => 
                           n6011);
   U5605 : AO7 port map( A => n6024, B => n5918, C => n6025, Z => n6023);
   U5606 : AO3 port map( A => n5863, B => n5929, C => n6026, D => n4363, Z => 
                           n6022);
   U5607 : AO1 port map( A => n4831, B => n4801, C => n6027, D => n6028, Z => 
                           n6009);
   U5608 : AN3 port map( A => n5857, B => n5885, C => n5905, Z => n6028);
   U5609 : NR2 port map( A => n4358, B => n5932, Z => n6027);
   U5610 : IV port map( A => n6029, Z => n5975);
   U5611 : AO7 port map( A => n6030, B => n5009, C => n6031, Z => n4173);
   U5612 : AO2 port map( A => n5823, B => n4693, C => n7807, D => n5824, Z => 
                           n6031);
   U5613 : MUX21L port map( A => n6032, B => n6033, S => n4395, Z => n4693);
   U5614 : AO1 port map( A => n6034, B => n6035, C => n6036, D => n6037, Z => 
                           n6033);
   U5615 : AO1 port map( A => n5895, B => n4801, C => n6038, D => n6039, Z => 
                           n6037);
   U5616 : AO4 port map( A => n5929, B => n6008, C => n6040, D => n4805, Z => 
                           n6039);
   U5617 : AO7 port map( A => n5918, B => n4832, C => n5842, Z => n6038);
   U5618 : IV port map( A => n5990, Z => n4832);
   U5619 : AO4 port map( A => n6041, B => n5852, C => n6042, D => n5858, Z => 
                           n6036);
   U5620 : AO1 port map( A => n5873, B => n6043, C => n6044, D => n6045, Z => 
                           n6042);
   U5621 : AN3 port map( A => n5925, B => n5885, C => n6046, Z => n6045);
   U5622 : AO4 port map( A => n5921, B => n6047, C => n5929, D => n6048, Z => 
                           n6044);
   U5623 : ND2 port map( A => n6002, B => n5866, Z => n6043);
   U5624 : AO1 port map( A => n5873, B => n5919, C => n6049, D => n6050, Z => 
                           n6041);
   U5625 : AO6 port map( A => n5974, B => n6046, C => n5929, Z => n6050);
   U5626 : AO4 port map( A => n4805, B => n5933, C => n5921, D => n5861, Z => 
                           n6049);
   U5627 : IV port map( A => n6051, Z => n5919);
   U5628 : AO1 port map( A => n5857, B => n6052, C => n6001, D => n5936, Z => 
                           n6035);
   U5629 : NR2 port map( A => n5836, B => n5921, Z => n5936);
   U5630 : NR2 port map( A => n5883, B => n5921, Z => n6001);
   U5631 : ND2 port map( A => n4806, B => n6053, Z => n6052);
   U5632 : AO1 port map( A => n6018, B => n5873, C => n4808, D => n6054, Z => 
                           n6034);
   U5633 : AO6 port map( A => n5944, B => n6008, C => n4805, Z => n6054);
   U5634 : AO1 port map( A => n4820, B => n6055, C => n6056, D => n6057, Z => 
                           n6032);
   U5635 : AO4 port map( A => n6058, B => n4800, C => n6059, D => n5852, Z => 
                           n6057);
   U5636 : IV port map( A => n6060, Z => n5852);
   U5637 : AO1 port map( A => n5873, B => n5955, C => n6061, D => n5996, Z => 
                           n6059);
   U5638 : NR2 port map( A => n5955, B => n4805, Z => n5996);
   U5639 : AO4 port map( A => v_RAM_OUT0_18_port, B => n5836, C => n5921, D => 
                           n6019, Z => n6061);
   U5640 : IV port map( A => n6062, Z => n5955);
   U5641 : AO1 port map( A => n6000, B => n4358, C => n6063, D => n6064, Z => 
                           n6058);
   U5642 : AN3 port map( A => n5942, B => n5932, C => n5925, Z => n6064);
   U5643 : NR2 port map( A => v_RAM_OUT0_20_port, B => n5944, Z => n6063);
   U5644 : ND4 port map( A => n6065, B => n6066, C => n6067, D => n4797, Z => 
                           n6056);
   U5645 : ND4 port map( A => n5857, B => n6068, C => n5836, D => n4403, Z => 
                           n6067);
   U5646 : IV port map( A => n5868, Z => n5836);
   U5647 : ND3 port map( A => n6002, B => n5883, C => n5846, Z => n6066);
   U5648 : AO7 port map( A => n6069, B => n5884, C => n4804, Z => n6065);
   U5649 : NR3 port map( A => n4808, B => n4409, C => n5905, Z => n6069);
   U5650 : IV port map( A => n6070, Z => n5905);
   U5651 : AO3 port map( A => n5918, B => n6071, C => n6072, D => n6073, Z => 
                           n6055);
   U5652 : AO2 port map( A => n4801, B => n6074, C => n6075, D => n5857, Z => 
                           n6073);
   U5653 : ND2 port map( A => n5989, B => n5958, Z => n6074);
   U5654 : ND3 port map( A => n5859, B => n5974, C => n5925, Z => n6072);
   U5655 : ND2 port map( A => n5942, B => n5932, Z => n6071);
   U5656 : AO7 port map( A => n6076, B => n5009, C => n6077, Z => n4172);
   U5657 : AO2 port map( A => n5823, B => n4696, C => n7865, D => n5824, Z => 
                           n6077);
   U5658 : IV port map( A => n6078, Z => n4696);
   U5659 : AO7 port map( A => n6079, B => n5827, C => n6080, Z => n6078);
   U5660 : MUX21L port map( A => n6081, B => n6082, S => n4395, Z => n6080);
   U5661 : ND4 port map( A => n6083, B => n6084, C => n6085, D => n6086, Z => 
                           n6082);
   U5662 : AO2 port map( A => n4794, B => n6087, C => n6088, D => n6089, Z => 
                           n6086);
   U5663 : ND2 port map( A => n6019, B => n6008, Z => n6087);
   U5664 : IV port map( A => n6090, Z => n6085);
   U5665 : AO4 port map( A => n6091, B => n5942, C => n5954, D => n6092, Z => 
                           n6090);
   U5666 : EO1 port map( A => n5994, B => n5987, C => n4797, D => n5970, Z => 
                           n6084);
   U5667 : NR2 port map( A => n5973, B => n5882, Z => n5970);
   U5668 : ND2 port map( A => n5974, B => n6068, Z => n5987);
   U5669 : AO2 port map( A => n5846, B => n6093, C => n5884, D => n5856, Z => 
                           n6083);
   U5670 : NR4 port map( A => n6094, B => n6095, C => n6096, D => n6097, Z => 
                           n6081);
   U5671 : AO4 port map( A => n6098, B => n6099, C => n5832, D => n5962, Z => 
                           n6097);
   U5672 : AO3 port map( A => n6100, B => n5963, C => v_RAM_OUT0_21_port, D => 
                           n6101, Z => n6099);
   U5673 : EO1 port map( A => n6102, B => n5861, C => n5898, D => n6103, Z => 
                           n6101);
   U5674 : IV port map( A => n5841, Z => n5861);
   U5675 : NR2 port map( A => n4802, B => n5881, Z => n5841);
   U5676 : AO3 port map( A => n6104, B => n5892, C => n6105, D => n6106, Z => 
                           n6098);
   U5677 : AO2 port map( A => n5961, B => n6107, C => n6108, D => n6109, Z => 
                           n6106);
   U5678 : ND2 port map( A => n6002, B => n6047, Z => n6109);
   U5679 : ND2 port map( A => n4804, B => n5995, Z => n6107);
   U5680 : AO2 port map( A => n6110, B => n5951, C => n6111, D => n6112, Z => 
                           n6105);
   U5681 : NR2 port map( A => n4822, B => n5973, Z => n6110);
   U5682 : NR2 port map( A => n6113, B => n5869, Z => n6104);
   U5683 : AO4 port map( A => n5856, B => n5839, C => n5922, D => n5983, Z => 
                           n6096);
   U5684 : AO4 port map( A => n5862, B => n5870, C => n6092, D => n6114, Z => 
                           n6095);
   U5685 : AO3 port map( A => n5939, B => n6091, C => n6115, D => n6116, Z => 
                           n6094);
   U5686 : ND3 port map( A => n5989, B => n5958, C => n6089, Z => n6116);
   U5687 : OR3 port map( A => n6088, B => n5956, C => n4797, Z => n6115);
   U5688 : AO1 port map( A => n6117, B => n4804, C => n6118, D => n6119, Z => 
                           n6079);
   U5689 : AO4 port map( A => n6120, B => n6121, C => n5890, D => n5902, Z => 
                           n6119);
   U5690 : ND2 port map( A => n6047, B => n5855, Z => n5902);
   U5691 : AO6 port map( A => n5972, B => n6122, C => n5951, Z => n6120);
   U5692 : NR2 port map( A => n4363, B => v_RAM_OUT0_18_port, Z => n5972);
   U5693 : AO7 port map( A => n5901, B => n5883, C => n6123, Z => n6118);
   U5694 : AO2 port map( A => n5969, B => n6122, C => n6102, D => n6124, Z => 
                           n6123);
   U5695 : ND2 port map( A => n4806, B => n5942, Z => n6122);
   U5696 : AO7 port map( A => n5879, B => n5898, C => n5892, Z => n6117);
   U5697 : AO7 port map( A => n6125, B => n5009, C => n6126, Z => n4171);
   U5698 : AO2 port map( A => n5823, B => n4699, C => n7874, D => n5824, Z => 
                           n6126);
   U5699 : MUX21L port map( A => n6127, B => n4792, S => n4395, Z => n4699);
   U5700 : ND4 port map( A => n6128, B => n6129, C => n6130, D => n6131, Z => 
                           n4792);
   U5701 : AO1 port map( A => n6060, B => n6132, C => n6133, D => n6134, Z => 
                           n6131);
   U5702 : AO4 port map( A => n6135, B => n5858, C => n6103, D => n4797, Z => 
                           n6134);
   U5703 : NR2 port map( A => n6136, B => n5869, Z => n6103);
   U5704 : IV port map( A => n4820, Z => n5858);
   U5705 : NR2 port map( A => n6137, B => n6138, Z => n6135);
   U5706 : AO4 port map( A => n6020, B => n5921, C => n5918, D => n6021, Z => 
                           n6138);
   U5707 : ND2 port map( A => n6100, B => n6008, Z => n6021);
   U5708 : EON1 port map( A => n6040, B => n4805, C => n6139, D => n5857, Z => 
                           n6137);
   U5709 : NR2 port map( A => n5881, B => n6088, Z => n6040);
   U5710 : AO4 port map( A => n5832, B => n6019, C => n5839, D => n5958, Z => 
                           n6133);
   U5711 : IV port map( A => n6140, Z => n5958);
   U5712 : IV port map( A => n4794, Z => n5839);
   U5713 : AO3 port map( A => n4805, B => n6046, C => n6025, D => n6141, Z => 
                           n6132);
   U5714 : AO2 port map( A => n5857, B => n6142, C => n5873, D => n6143, Z => 
                           n6141);
   U5715 : ND2 port map( A => n6008, B => n6005, Z => n6143);
   U5716 : ND2 port map( A => n5974, B => n5866, Z => n6142);
   U5717 : IV port map( A => n5928, Z => n5866);
   U5718 : AO2 port map( A => n5925, B => n5956, C => n5954, D => n4801, Z => 
                           n6025);
   U5719 : ND2 port map( A => n6046, B => n5867, Z => n5954);
   U5720 : AO2 port map( A => n6089, B => n6018, C => n6144, D => n5922, Z => 
                           n6130);
   U5721 : AO7 port map( A => n5994, B => n4794, C => n6145, Z => n6129);
   U5722 : AO2 port map( A => n6146, B => n5846, C => n5845, D => n6147, Z => 
                           n6128);
   U5723 : ND2 port map( A => n5832, B => n6092, Z => n6147);
   U5724 : NR2 port map( A => n5959, B => n6070, Z => n6146);
   U5725 : AO3 port map( A => n6148, B => n4797, C => n6149, D => n6150, Z => 
                           n6127);
   U5726 : AO2 port map( A => n5844, B => n4809, C => v_RAM_OUT0_21_port, D => 
                           n4807, Z => n6150);
   U5727 : ND4 port map( A => n6151, B => n6152, C => n6153, D => n6154, Z => 
                           n4807);
   U5728 : AO2 port map( A => n6155, B => n6102, C => n6108, D => n6156, Z => 
                           n6154);
   U5729 : ND2 port map( A => n5885, B => n6005, Z => n6156);
   U5730 : IV port map( A => n6088, Z => n6005);
   U5731 : NR2 port map( A => n4367, B => v_RAM_OUT0_16_port, Z => n6088);
   U5732 : NR2 port map( A => n6140, B => n4793, Z => n6155);
   U5733 : AO2 port map( A => n5957, B => n6157, C => n6112, D => n5915, Z => 
                           n6153);
   U5734 : ND2 port map( A => n5942, B => n5931, Z => n5915);
   U5735 : AO2 port map( A => n5951, B => n5885, C => n5960, D => n6019, Z => 
                           n6152);
   U5736 : AO2 port map( A => n5969, B => n5856, C => n5961, D => n5962, Z => 
                           n6151);
   U5737 : AO3 port map( A => n4830, B => n4804, C => n6158, D => n6159, Z => 
                           n4809);
   U5738 : AO2 port map( A => n5928, B => n5925, C => n6160, D => n4801, Z => 
                           n6159);
   U5739 : NR2 port map( A => n5995, B => v_RAM_OUT0_16_port, Z => n5928);
   U5740 : ND2 port map( A => n5857, B => n5944, Z => n6158);
   U5741 : AO2 port map( A => n4794, B => n6161, C => n5842, D => n6162, Z => 
                           n6149);
   U5742 : AO3 port map( A => n5921, B => n4802, C => n6163, D => n6026, Z => 
                           n6162);
   U5743 : IV port map( A => n5940, Z => n6026);
   U5744 : NR2 port map( A => n6047, B => n4805, Z => n5940);
   U5745 : ND2 port map( A => n5938, B => n5925, Z => n6163);
   U5746 : ND2 port map( A => n5855, B => n6068, Z => n6161);
   U5747 : IV port map( A => n5891, Z => n6068);
   U5748 : IV port map( A => n5938, Z => n5855);
   U5749 : AO7 port map( A => n6164, B => n5009, C => n6165, Z => n4170);
   U5750 : AO2 port map( A => n5823, B => n4702, C => n7873, D => n5824, Z => 
                           n6165);
   U5751 : IV port map( A => n6166, Z => n4702);
   U5752 : AO7 port map( A => n6167, B => n5827, C => n6168, Z => n6166);
   U5753 : MUX21L port map( A => n6169, B => n6170, S => n4395, Z => n6168);
   U5754 : ND4 port map( A => n6171, B => n6172, C => n6173, D => n6174, Z => 
                           n6170);
   U5755 : AO2 port map( A => n6111, B => n6144, C => n5994, D => n6175, Z => 
                           n6174);
   U5756 : ND2 port map( A => n6100, B => n5933, Z => n6175);
   U5757 : NR2 port map( A => n5939, B => n6136, Z => n6111);
   U5758 : AO2 port map( A => n5846, B => n6176, C => n6089, D => n5990, Z => 
                           n6173);
   U5759 : NR2 port map( A => n4800, B => n4805, Z => n6089);
   U5760 : ND2 port map( A => n6002, B => n5856, Z => n6176);
   U5761 : IV port map( A => n5869, Z => n5856);
   U5762 : EO1 port map( A => n5835, B => n6114, C => n5832, D => n5863, Z => 
                           n6172);
   U5763 : NR2 port map( A => n5869, B => n6140, Z => n5863);
   U5764 : ND2 port map( A => n6019, B => n6053, Z => n6114);
   U5765 : IV port map( A => n6113, Z => n6053);
   U5766 : AO2 port map( A => n6177, B => n6019, C => n4794, D => n6093, Z => 
                           n6171);
   U5767 : IV port map( A => n5895, Z => n6093);
   U5768 : NR4 port map( A => n6178, B => n6179, C => n6180, D => n6181, Z => 
                           n6169);
   U5769 : AO4 port map( A => n6182, B => n6183, C => n5832, D => n6000, Z => 
                           n6181);
   U5770 : OR2 port map( A => n6018, B => n6140, Z => n6000);
   U5771 : AO3 port map( A => n5898, B => n6184, C => v_RAM_OUT0_21_port, D => 
                           n6185, Z => n6183);
   U5772 : AO2 port map( A => n5961, B => n4798, C => n5960, D => n5944, Z => 
                           n6185);
   U5773 : IV port map( A => n6148, Z => n4798);
   U5774 : NR2 port map( A => n4802, B => n5956, Z => n6148);
   U5775 : AO3 port map( A => n5894, B => n5933, C => n6186, D => n6187, Z => 
                           n6182);
   U5776 : EO1 port map( A => n6102, B => v_RAM_OUT0_19_port, C => n5883, D => 
                           n5903, Z => n6187);
   U5777 : EO1 port map( A => n6188, B => n6108, C => n5963, D => n5897, Z => 
                           n6186);
   U5778 : NR2 port map( A => n6018, B => n5868, Z => n5897);
   U5779 : IV port map( A => n5969, Z => n5963);
   U5780 : NR2 port map( A => n5922, B => n6136, Z => n6188);
   U5781 : MUX21L port map( A => n6091, B => n6189, S => n5870, Z => n6180);
   U5782 : NR2 port map( A => n6190, B => n4794, Z => n6189);
   U5783 : NR2 port map( A => n4800, B => n5918, Z => n4794);
   U5784 : AN3 port map( A => n4793, B => v_RAM_OUT0_18_port, C => n5842, Z => 
                           n6190);
   U5785 : IV port map( A => n6144, Z => n6091);
   U5786 : NR2 port map( A => n4808, B => n4805, Z => n6144);
   U5787 : AO4 port map( A => n5983, B => n5843, C => n6075, D => n5862, Z => 
                           n6179);
   U5788 : IV port map( A => n5994, Z => n5862);
   U5789 : NR2 port map( A => n4808, B => n5929, Z => n5994);
   U5790 : NR2 port map( A => n5879, B => n6140, Z => n6075);
   U5791 : NR2 port map( A => n4802, B => n4354, Z => n6140);
   U5792 : ND2 port map( A => n5906, B => n5989, Z => n5843);
   U5793 : IV port map( A => n5846, Z => n5983);
   U5794 : AO4 port map( A => n6092, B => n4806, C => n4797, D => n6191, Z => 
                           n6178);
   U5795 : ND2 port map( A => n5974, B => n5859, Z => n6191);
   U5796 : IV port map( A => n6160, Z => n5859);
   U5797 : IV port map( A => n5845, Z => n5974);
   U5798 : IV port map( A => n6177, Z => n4797);
   U5799 : NR2 port map( A => n4800, B => n5929, Z => n6177);
   U5800 : IV port map( A => n5835, Z => n6092);
   U5801 : NR2 port map( A => n4800, B => n5921, Z => n5835);
   U5802 : IV port map( A => n5842, Z => n4800);
   U5803 : ND2 port map( A => v_RAM_OUT0_21_port, B => n4395, Z => n5827);
   U5804 : NR4 port map( A => n6192, B => n6193, C => n6194, D => n6195, Z => 
                           n6167);
   U5805 : AO4 port map( A => n5896, B => n6048, C => n5895, D => n5894, Z => 
                           n6195);
   U5806 : IV port map( A => n5951, Z => n5894);
   U5807 : NR2 port map( A => n6113, B => n6070, Z => n5895);
   U5808 : NR2 port map( A => v_RAM_OUT0_16_port, B => n5880, Z => n6070);
   U5809 : IV port map( A => n4831, Z => n6048);
   U5810 : IV port map( A => n6102, Z => n5896);
   U5811 : EON1 port map( A => n5890, B => n6157, C => n5876, D => n5969, Z => 
                           n6194);
   U5812 : IV port map( A => n5961, Z => n5890);
   U5813 : EON1 port map( A => n6196, B => n5898, C => n6006, D => n6112, Z => 
                           n6193);
   U5814 : ND2 port map( A => n5989, B => n5867, Z => n6006);
   U5815 : IV port map( A => n4793, Z => n5989);
   U5816 : IV port map( A => n5957, Z => n5898);
   U5817 : NR2 port map( A => n5869, B => n4822, Z => n6196);
   U5818 : AO4 port map( A => n6197, B => n5892, C => n5901, D => n6198, Z => 
                           n6192);
   U5819 : ND2 port map( A => n6008, B => n5944, Z => n6198);
   U5820 : IV port map( A => n5956, Z => n6008);
   U5821 : NR2 port map( A => n4354, B => n5880, Z => n5956);
   U5822 : IV port map( A => n6108, Z => n5901);
   U5823 : NR2 port map( A => n6160, B => n5831, Z => n6197);
   U5824 : NR2 port map( A => n6100, B => v_RAM_OUT0_16_port, Z => n6160);
   U5825 : AO7 port map( A => n6199, B => n5009, C => n6200, Z => n4169);
   U5826 : AO2 port map( A => n5823, B => n4705, C => n7806, D => n5824, Z => 
                           n6200);
   U5827 : MUX21L port map( A => n6201, B => n6202, S => n4395, Z => n4705);
   U5828 : AO6 port map( A => v_RAM_OUT0_21_port, B => n6203, C => n4818, Z => 
                           n6202);
   U5829 : AO3 port map( A => n5870, B => n6204, C => n6205, D => n6206, Z => 
                           n4818);
   U5830 : ND4 port map( A => n6207, B => n6208, C => n6209, D => n6210, Z => 
                           n6206);
   U5831 : NR2 port map( A => v_RAM_OUT0_21_port, B => n6211, Z => n6210);
   U5832 : AO6 port map( A => n5885, B => n6046, C => n5929, Z => n6211);
   U5833 : IV port map( A => n5973, Z => n6046);
   U5834 : NR2 port map( A => v_RAM_OUT0_16_port, B => n5879, Z => n5973);
   U5835 : IV port map( A => n4822, Z => n5885);
   U5836 : AO2 port map( A => n6112, B => n6139, C => n5960, D => n6157, Z => 
                           n6209);
   U5837 : ND2 port map( A => n6047, B => n5933, Z => n6157);
   U5838 : IV port map( A => n5881, Z => n5933);
   U5839 : NR2 port map( A => n4354, B => n5879, Z => n5881);
   U5840 : ND2 port map( A => n4804, B => n6047, Z => n6139);
   U5841 : IV port map( A => n6136, Z => n4804);
   U5842 : AO2 port map( A => n6113, B => n5961, C => n6102, D => n5879, Z => 
                           n6208);
   U5843 : NR2 port map( A => n4354, B => n4412, Z => n6113);
   U5844 : AO2 port map( A => n6108, B => n5942, C => n5969, D => n4367, Z => 
                           n6207);
   U5845 : ND3 port map( A => n6060, B => n6212, C => n6213, Z => n6205);
   U5846 : AO1 port map( A => n4822, B => n5857, C => n5869, D => n6214, Z => 
                           n6213);
   U5847 : NR2 port map( A => n5938, B => n5918, Z => n6214);
   U5848 : NR2 port map( A => n6100, B => n4354, Z => n5938);
   U5849 : IV port map( A => n6124, Z => n6100);
   U5850 : NR2 port map( A => v_RAM_OUT0_19_port, B => v_RAM_OUT0_16_port, Z =>
                           n5869);
   U5851 : AO4 port map( A => n5845, B => n5893, C => n4801, D => n6215, Z => 
                           n6212);
   U5852 : NR2 port map( A => v_RAM_OUT0_20_port, B => n6019, Z => n6215);
   U5853 : IV port map( A => n5893, Z => n6019);
   U5854 : NR2 port map( A => v_RAM_OUT0_16_port, B => n6124, Z => n5893);
   U5855 : NR2 port map( A => n4403, B => v_RAM_OUT0_17_port, Z => n6060);
   U5856 : ND2 port map( A => n4820, B => n4830, Z => n6204);
   U5857 : IV port map( A => n4819, Z => n4830);
   U5858 : NR2 port map( A => n4363, B => n4403, Z => n4820);
   U5859 : IV port map( A => n6216, Z => n5870);
   U5860 : AO4 port map( A => n4822, B => n5892, C => n5903, D => n4823, Z => 
                           n6203);
   U5861 : IV port map( A => n6024, Z => n4823);
   U5862 : NR2 port map( A => n5831, B => n5891, Z => n6024);
   U5863 : NR2 port map( A => n4802, B => v_RAM_OUT0_16_port, Z => n5891);
   U5864 : IV port map( A => n6112, Z => n5903);
   U5865 : IV port map( A => n5960, Z => n5892);
   U5866 : NR2 port map( A => n5918, B => n4363, Z => n5960);
   U5867 : AO3 port map( A => n5990, B => n5832, C => n6217, D => n6218, Z => 
                           n6201);
   U5868 : AO2 port map( A => n5842, B => n4826, C => v_RAM_OUT0_21_port, D => 
                           n4833, Z => n6218);
   U5869 : ND4 port map( A => n6219, B => n6220, C => n6221, D => n6222, Z => 
                           n4833);
   U5870 : AO2 port map( A => v_RAM_OUT0_17_port, B => n6223, C => n6051, D => 
                           n6102, Z => n6222);
   U5871 : NR2 port map( A => n4805, B => v_RAM_OUT0_17_port, Z => n6102);
   U5872 : AO4 port map( A => n4409, B => n5883, C => n6224, D => n4358, Z => 
                           n6223);
   U5873 : NR2 port map( A => n5900, B => n5959, Z => n6224);
   U5874 : ND2 port map( A => n4354, B => n5932, Z => n5883);
   U5875 : AO2 port map( A => n5957, B => n5876, C => n5951, D => n6184, Z => 
                           n6221);
   U5876 : IV port map( A => n6020, Z => n6184);
   U5877 : NR2 port map( A => n5882, B => n6145, Z => n6020);
   U5878 : NR2 port map( A => n5929, B => n4363, Z => n5951);
   U5879 : ND2 port map( A => n6047, B => n5906, Z => n5876);
   U5880 : IV port map( A => n5959, Z => n5906);
   U5881 : NR2 port map( A => n4354, B => n5995, Z => n5959);
   U5882 : IV port map( A => n5880, Z => n5995);
   U5883 : NR2 port map( A => n5929, B => v_RAM_OUT0_17_port, Z => n5957);
   U5884 : AO2 port map( A => n6112, B => n5942, C => n6136, D => n5961, Z => 
                           n6220);
   U5885 : NR2 port map( A => n4805, B => n4363, Z => n5961);
   U5886 : IV port map( A => n5925, Z => n4805);
   U5887 : NR2 port map( A => n4354, B => n6124, Z => n6136);
   U5888 : ND2 port map( A => v_RAM_OUT0_16_port, B => n4802, Z => n5942);
   U5889 : IV port map( A => n5922, Z => n4802);
   U5890 : NR2 port map( A => n4363, B => n5921, Z => n6112);
   U5891 : AO2 port map( A => n5969, B => n5922, C => n6108, D => n5962, Z => 
                           n6219);
   U5892 : ND2 port map( A => n6002, B => n4806, Z => n5962);
   U5893 : IV port map( A => n6145, Z => n4806);
   U5894 : NR2 port map( A => v_RAM_OUT0_22_port, B => v_RAM_OUT0_16_port, Z =>
                           n6145);
   U5895 : IV port map( A => n5831, Z => n6002);
   U5896 : NR2 port map( A => n5932, B => n4354, Z => n5831);
   U5897 : NR2 port map( A => n5921, B => v_RAM_OUT0_17_port, Z => n6108);
   U5898 : NR2 port map( A => n5918, B => v_RAM_OUT0_17_port, Z => n5969);
   U5899 : AO7 port map( A => n6062, B => n5929, C => n6225, Z => n4826);
   U5900 : AO2 port map( A => n6216, B => n6226, C => n6051, D => n4801, Z => 
                           n6225);
   U5901 : NR2 port map( A => n4822, B => n6124, Z => n6051);
   U5902 : AO7 port map( A => n4358, B => n5931, C => n5918, Z => n6226);
   U5903 : IV port map( A => n5900, Z => n5931);
   U5904 : NR2 port map( A => n5944, B => v_RAM_OUT0_16_port, Z => n5900);
   U5905 : IV port map( A => n5879, Z => n5944);
   U5906 : NR2 port map( A => n5845, B => n4793, Z => n6216);
   U5907 : NR2 port map( A => n4354, B => v_RAM_OUT0_19_port, Z => n5845);
   U5908 : IV port map( A => n5857, Z => n5929);
   U5909 : NR2 port map( A => n5882, B => n6018, Z => n6062);
   U5910 : NR2 port map( A => n5932, B => v_RAM_OUT0_16_port, Z => n6018);
   U5911 : IV port map( A => n5939, Z => n5932);
   U5912 : NR2 port map( A => n4367, B => n4354, Z => n5882);
   U5913 : NR2 port map( A => v_RAM_OUT0_21_port, B => v_RAM_OUT0_17_port, Z =>
                           n5842);
   U5914 : AO2 port map( A => n6227, B => n5844, C => n4831, D => n5846, Z => 
                           n6217);
   U5915 : NR2 port map( A => n4808, B => n5918, Z => n5846);
   U5916 : IV port map( A => n5873, Z => n5918);
   U5917 : NR2 port map( A => n4358, B => v_RAM_OUT0_20_port, Z => n5873);
   U5918 : NR2 port map( A => n5880, B => n4822, Z => n4831);
   U5919 : NR2 port map( A => n4354, B => n5939, Z => n4822);
   U5920 : NR2 port map( A => n4412, B => v_RAM_OUT0_19_port, Z => n5880);
   U5921 : NR2 port map( A => n4829, B => n4819, Z => n6227);
   U5922 : NR2 port map( A => n5925, B => n5857, Z => n4819);
   U5923 : NR2 port map( A => v_RAM_OUT0_20_port, B => v_RAM_OUT0_18_port, Z =>
                           n5857);
   U5924 : NR2 port map( A => n4358, B => n4409, Z => n5925);
   U5925 : IV port map( A => n6121, Z => n4829);
   U5926 : ND2 port map( A => n6047, B => n5867, Z => n6121);
   U5927 : ND2 port map( A => n5879, B => v_RAM_OUT0_16_port, Z => n5867);
   U5928 : NR2 port map( A => n4367, B => v_RAM_OUT0_22_port, Z => n5879);
   U5929 : ND2 port map( A => v_RAM_OUT0_22_port, B => n4354, Z => n6047);
   U5930 : IV port map( A => n5884, Z => n5832);
   U5931 : NR2 port map( A => n4808, B => n5921, Z => n5884);
   U5932 : IV port map( A => n4801, Z => n5921);
   U5933 : NR2 port map( A => n4409, B => v_RAM_OUT0_18_port, Z => n4801);
   U5934 : IV port map( A => n5844, Z => n4808);
   U5935 : NR2 port map( A => n4363, B => v_RAM_OUT0_21_port, Z => n5844);
   U5936 : NR2 port map( A => n4793, B => n5868, Z => n5990);
   U5937 : NR2 port map( A => n4354, B => v_RAM_OUT0_22_port, Z => n5868);
   U5938 : NR2 port map( A => v_RAM_OUT0_16_port, B => n5922, Z => n4793);
   U5939 : NR2 port map( A => n5939, B => n6124, Z => n5922);
   U5940 : NR2 port map( A => n4367, B => n4412, Z => n6124);
   U5941 : NR2 port map( A => v_RAM_OUT0_22_port, B => v_RAM_OUT0_19_port, Z =>
                           n5939);
   U5942 : NR2 port map( A => n5384, B => n5824, Z => n5823);
   U5943 : NR2 port map( A => n5384, B => n4733, Z => n5824);
   U5944 : AN3 port map( A => n4560, B => v_CALCULATION_CNTR_0_port, C => n6228
                           , Z => n4733);
   U5945 : AO7 port map( A => n6229, B => n5009, C => n6230, Z => n4168);
   U5946 : AO2 port map( A => n6231, B => n4709, C => n7900, D => n6232, Z => 
                           n6230);
   U5947 : IV port map( A => n6233, Z => n4709);
   U5948 : AO7 port map( A => n6234, B => n6235, C => n6236, Z => n6233);
   U5949 : MUX21L port map( A => n6237, B => n6238, S => n4396, Z => n6236);
   U5950 : AO3 port map( A => n6239, B => n6240, C => n6241, D => n6242, Z => 
                           n6238);
   U5951 : AO1 port map( A => n6243, B => n6244, C => n6245, D => n6246, Z => 
                           n6242);
   U5952 : AO6 port map( A => n6247, B => n6248, C => n6249, Z => n6246);
   U5953 : ND3 port map( A => v_RAM_OUT0_26_port, B => n6250, C => n6239, Z => 
                           n6248);
   U5954 : AN3 port map( A => n6251, B => n4359, C => n6252, Z => n6245);
   U5955 : EO1 port map( A => n6253, B => n6254, C => n4971, D => n6255, Z => 
                           n6241);
   U5956 : NR4 port map( A => n6256, B => n6257, C => n6258, D => n6259, Z => 
                           n6237);
   U5957 : AO4 port map( A => n6260, B => n6261, C => n4971, D => n6262, Z => 
                           n6259);
   U5958 : ND2 port map( A => n6263, B => n6264, Z => n6262);
   U5959 : ND2 port map( A => n6265, B => n4980, Z => n6261);
   U5960 : NR3 port map( A => n6266, B => v_RAM_OUT0_28_port, C => n6267, Z => 
                           n6258);
   U5961 : AO4 port map( A => n6268, B => n4979, C => n6269, D => n6270, Z => 
                           n6257);
   U5962 : AO1 port map( A => n6271, B => n6252, C => n6272, D => n6273, Z => 
                           n6268);
   U5963 : AO6 port map( A => n6274, B => n6275, C => n6266, Z => n6273);
   U5964 : AO4 port map( A => n6249, B => n4974, C => n6255, D => n6260, Z => 
                           n6272);
   U5965 : NR2 port map( A => n6276, B => n6277, Z => n6255);
   U5966 : AO3 port map( A => n6278, B => n6247, C => n6279, D => n6280, Z => 
                           n6256);
   U5967 : AO2 port map( A => n6281, B => n6282, C => n4975, D => n6283, Z => 
                           n6280);
   U5968 : AO3 port map( A => n4974, B => n6284, C => n6285, D => n6286, Z => 
                           n6283);
   U5969 : ND2 port map( A => n4994, B => n6287, Z => n6286);
   U5970 : OR3 port map( A => n6288, B => n6289, C => n6260, Z => n6285);
   U5971 : AO4 port map( A => n6290, B => n6266, C => n6260, D => n6291, Z => 
                           n6282);
   U5972 : MUX21L port map( A => n6292, B => n6254, S => n6293, Z => n6279);
   U5973 : NR4 port map( A => n6294, B => n6295, C => n6296, D => n6297, Z => 
                           n6234);
   U5974 : AO4 port map( A => n6298, B => n6264, C => n6299, D => n6300, Z => 
                           n6297);
   U5975 : AO4 port map( A => n6301, B => n6302, C => n6303, D => n6304, Z => 
                           n6296);
   U5976 : AO4 port map( A => n6305, B => n6306, C => n4359, D => n6307, Z => 
                           n6295);
   U5977 : MUX21L port map( A => n4996, B => n6308, S => n4364, Z => n6307);
   U5978 : AO4 port map( A => n6309, B => n6310, C => n6311, D => n6312, Z => 
                           n6294);
   U5979 : ND2 port map( A => n6313, B => n6314, Z => n6312);
   U5980 : AO7 port map( A => n6315, B => n5009, C => n6316, Z => n4167);
   U5981 : AO2 port map( A => n6231, B => n4714, C => n7906, D => n6232, Z => 
                           n6316);
   U5982 : MUX21L port map( A => n6317, B => n6318, S => n4396, Z => n4714);
   U5983 : AO1 port map( A => n6319, B => n6320, C => n6321, D => n6322, Z => 
                           n6318);
   U5984 : AO1 port map( A => n6265, B => n6323, C => n6324, D => n6325, Z => 
                           n6322);
   U5985 : AO4 port map( A => n6326, B => n6327, C => n6328, D => n6329, Z => 
                           n6325);
   U5986 : NR2 port map( A => n6290, B => n6308, Z => n6328);
   U5987 : AO7 port map( A => n6330, B => n4979, C => n6250, Z => n6324);
   U5988 : AO4 port map( A => n6331, B => n6266, C => n6332, D => n6260, Z => 
                           n6321);
   U5989 : AO1 port map( A => n6333, B => n4997, C => n6334, D => n6335, Z => 
                           n6332);
   U5990 : NR2 port map( A => v_RAM_OUT0_28_port, B => n6244, Z => n6335);
   U5991 : AO3 port map( A => n6336, B => n6337, C => n6338, D => n6339, Z => 
                           n6334);
   U5992 : ND3 port map( A => n6340, B => n6341, C => n4975, Z => n6338);
   U5993 : AO1 port map( A => n6342, B => n6281, C => n6343, D => n6344, Z => 
                           n6331);
   U5994 : AO4 port map( A => n6337, B => n6267, C => n6345, D => n4979, Z => 
                           n6343);
   U5995 : NR2 port map( A => n6346, B => n6308, Z => n6345);
   U5996 : NR2 port map( A => n6347, B => n6289, Z => n6342);
   U5997 : AO1 port map( A => n6347, B => n4975, C => n6348, D => n6349, Z => 
                           n6320);
   U5998 : NR2 port map( A => n4979, B => n6350, Z => n6349);
   U5999 : NR2 port map( A => n4982, B => n6351, Z => n6319);
   U6000 : MUX21L port map( A => n6337, B => n6326, S => n6352, Z => n6351);
   U6001 : MUX21L port map( A => n6353, B => n6354, S => n4404, Z => n6317);
   U6002 : AN3 port map( A => n6355, B => n6356, C => n6357, Z => n6354);
   U6003 : AO1 port map( A => n6358, B => n6359, C => n6360, D => n6361, Z => 
                           n6357);
   U6004 : NR4 port map( A => v_RAM_OUT0_26_port, B => v_RAM_OUT0_25_port, C =>
                           n6330, D => n4996, Z => n6361);
   U6005 : AO4 port map( A => n6311, B => n6362, C => n6304, D => n6363, Z => 
                           n6360);
   U6006 : NR2 port map( A => n6287, B => n6364, Z => n6358);
   U6007 : AO2 port map( A => n6365, B => n6366, C => n6367, D => n6368, Z => 
                           n6356);
   U6008 : EO1 port map( A => n6369, B => n6278, C => n6370, D => n6371, Z => 
                           n6355);
   U6009 : NR4 port map( A => n6372, B => n6373, C => n6374, D => n6375, Z => 
                           n6353);
   U6010 : AO4 port map( A => n6309, B => n4972, C => v_RAM_OUT0_25_port, D => 
                           n6274, Z => n6375);
   U6011 : MUX21L port map( A => n6304, B => n6376, S => n6263, Z => n6374);
   U6012 : AO6 port map( A => n6368, B => n6264, C => n6377, Z => n6376);
   U6013 : AO4 port map( A => n6275, B => n6306, C => n6378, D => n6379, Z => 
                           n6373);
   U6014 : AO6 port map( A => n6380, B => n6381, C => n6359, Z => n6379);
   U6015 : AO6 port map( A => n6382, B => n6267, C => n6298, Z => n6372);
   U6016 : AO7 port map( A => n6383, B => n5009, C => n6384, Z => n4166);
   U6017 : AO2 port map( A => n6231, B => n4717, C => n7912, D => n6232, Z => 
                           n6384);
   U6018 : MUX21H port map( A => n6385, B => n6386, S => v_RAM_OUT0_31_port, Z 
                           => n4717);
   U6019 : AO1 port map( A => n6387, B => n6388, C => n6389, D => n6390, Z => 
                           n6386);
   U6020 : AO4 port map( A => n6264, B => n6391, C => n6392, D => n6260, Z => 
                           n6390);
   U6021 : AO1 port map( A => n6299, B => n4975, C => n6393, D => n6394, Z => 
                           n6392);
   U6022 : AO7 port map( A => n6326, B => n6395, C => n6396, Z => n6394);
   U6023 : IV port map( A => n6344, Z => n6396);
   U6024 : AO4 port map( A => n6337, B => n6397, C => n6398, D => n4979, Z => 
                           n6393);
   U6025 : AO3 port map( A => n6399, B => n6266, C => n6400, D => n6401, Z => 
                           n6389);
   U6026 : AO2 port map( A => n6402, B => n6403, C => n6404, D => n6252, Z => 
                           n6401);
   U6027 : AO7 port map( A => n6254, B => n6292, C => n6346, Z => n6400);
   U6028 : AO1 port map( A => n6281, B => n5006, C => n6405, D => n6406, Z => 
                           n6399);
   U6029 : IV port map( A => n6407, Z => n6406);
   U6030 : AO6 port map( A => n6408, B => n6265, C => n6409, Z => n6407);
   U6031 : AO4 port map( A => n6329, B => n6410, C => n4979, D => n6291, Z => 
                           n6405);
   U6032 : AO1 port map( A => n6281, B => n6411, C => n6409, D => n6412, Z => 
                           n6388);
   U6033 : AO6 port map( A => n6340, B => n4978, C => n4979, Z => n6412);
   U6034 : ND2 port map( A => n6244, B => n6413, Z => n6411);
   U6035 : AO1 port map( A => n6265, B => n6414, C => n4974, D => n6415, Z => 
                           n6387);
   U6036 : NR2 port map( A => n6329, B => n6416, Z => n6415);
   U6037 : AO7 port map( A => n6417, B => n6266, C => n6418, Z => n6385);
   U6038 : MUX21L port map( A => n6419, B => n6420, S => n4404, Z => n6418);
   U6039 : NR4 port map( A => n6421, B => n6422, C => n6423, D => n6424, Z => 
                           n6420);
   U6040 : AO4 port map( A => n6301, B => n6298, C => n6291, D => n6371, Z => 
                           n6424);
   U6041 : MUX21L port map( A => n6300, B => n6306, S => n5006, Z => n6423);
   U6042 : AO4 port map( A => n6309, B => n6425, C => n6426, D => n6311, Z => 
                           n6422);
   U6043 : ND2 port map( A => n6427, B => n6382, Z => n6425);
   U6044 : EON1 port map( A => n6428, B => n6304, C => n6429, D => n6380, Z => 
                           n6421);
   U6045 : AO4 port map( A => n6430, B => n6431, C => n6298, D => n6416, Z => 
                           n6419);
   U6046 : AO7 port map( A => n6432, B => n6326, C => n6433, Z => n6431);
   U6047 : AO3 port map( A => n6271, B => n6337, C => n6434, D => n4364, Z => 
                           n6430);
   U6048 : AO1 port map( A => n5005, B => n4975, C => n6435, D => n6436, Z => 
                           n6417);
   U6049 : AN3 port map( A => n6265, B => n6293, C => n6313, Z => n6436);
   U6050 : NR2 port map( A => n4359, B => n6340, Z => n6435);
   U6051 : AO3 port map( A => n6437, B => n4371, C => n6438, D => n6439, Z => 
                           n4165);
   U6052 : AO6 port map( A => n6440, B => n6441, C => n6442, Z => n6439);
   U6053 : AO4 port map( A => n6443, B => n6444, C => n6445, D => n6446, Z => 
                           n6442);
   U6054 : EO port map( A => n6447, B => n6448, Z => n6445);
   U6055 : EO port map( A => n6449, B => n6450, Z => n6448);
   U6056 : EN port map( A => n6451, B => n6452, Z => n6450);
   U6057 : EN port map( A => n4707, B => n6453, Z => n6447);
   U6058 : EO port map( A => n6454, B => n6455, Z => n6443);
   U6059 : EN port map( A => n6456, B => n6457, Z => n6455);
   U6060 : EO port map( A => n6458, B => n6459, Z => n6454);
   U6061 : EO port map( A => n6460, B => n6461, Z => n6459);
   U6062 : EO port map( A => v_KEY_COLUMN_24_port, B => v_DATA_COLUMN_24_port, 
                           Z => n6441);
   U6063 : AO2 port map( A => n6462, B => n6463, C => n6464, D => n6465, Z => 
                           n6438);
   U6064 : EO port map( A => n6466, B => n6467, Z => n6465);
   U6065 : EN port map( A => n6468, B => n6469, Z => n6467);
   U6066 : EO port map( A => n6470, B => n6471, Z => n6466);
   U6067 : EN port map( A => n6472, B => n6229, Z => n6471);
   U6068 : EO port map( A => n6473, B => n6474, Z => n6463);
   U6069 : EO port map( A => n6475, B => n6476, Z => n6474);
   U6070 : EO port map( A => n6477, B => n6478, Z => n6476);
   U6071 : EN port map( A => n4950, B => n6479, Z => n6473);
   U6072 : MUX21L port map( A => n4420, B => n4371, S => n6480, Z => n4164);
   U6073 : MUX21H port map( A => t_STATE_RAM0_1_24_port, B => v_RAM_IN0_24_port
                           , S => n6481, Z => n4163);
   U6074 : MUX21H port map( A => t_STATE_RAM0_2_24_port, B => v_RAM_IN0_24_port
                           , S => n6482, Z => n4162);
   U6075 : MUX21H port map( A => t_STATE_RAM0_3_24_port, B => v_RAM_IN0_24_port
                           , S => n4498, Z => n4161);
   U6076 : AO3 port map( A => n4420, B => n6483, C => n6484, D => n6485, Z => 
                           n4160);
   U6077 : AO2 port map( A => n6486, B => t_STATE_RAM0_3_24_port, C => 
                           v_RAM_OUT0_24_port, D => n4513, Z => n6485);
   U6078 : AO2 port map( A => n4564, B => t_STATE_RAM0_1_24_port, C => n4563, D
                           => t_STATE_RAM0_2_24_port, Z => n6484);
   U6079 : IV port map( A => n6487, Z => n4159);
   U6080 : AO6 port map( A => n6232, B => n7918, C => n6488, Z => n6487);
   U6081 : IV port map( A => n6489, Z => n6488);
   U6082 : AO2 port map( A => n6231, B => n4720, C => n5384, D => n6490, Z => 
                           n6489);
   U6083 : MUX21L port map( A => n6491, B => n6492, S => n4396, Z => n4720);
   U6084 : AO1 port map( A => n6493, B => n6494, C => n6495, D => n6496, Z => 
                           n6492);
   U6085 : AO1 port map( A => n6303, B => n4975, C => n6497, D => n6498, Z => 
                           n6496);
   U6086 : AO4 port map( A => n6337, B => n6416, C => n6499, D => n4979, Z => 
                           n6498);
   U6087 : AO7 port map( A => n6326, B => n5006, C => n6250, Z => n6497);
   U6088 : IV port map( A => n6398, Z => n5006);
   U6089 : AO4 port map( A => n6500, B => n6260, C => n6501, D => n6266, Z => 
                           n6495);
   U6090 : AO1 port map( A => n6281, B => n6502, C => n6503, D => n6504, Z => 
                           n6501);
   U6091 : AN3 port map( A => n6333, B => n6293, C => n6505, Z => n6504);
   U6092 : AO4 port map( A => n6329, B => n6506, C => n6337, D => n6507, Z => 
                           n6503);
   U6093 : ND2 port map( A => n6410, B => n6274, Z => n6502);
   U6094 : AO1 port map( A => n6281, B => n6327, C => n6508, D => n6509, Z => 
                           n6500);
   U6095 : AO6 port map( A => n6382, B => n6505, C => n6337, Z => n6509);
   U6096 : AO4 port map( A => n4979, B => n6341, C => n6329, D => n6269, Z => 
                           n6508);
   U6097 : IV port map( A => n6510, Z => n6327);
   U6098 : AO1 port map( A => n6265, B => n6511, C => n6409, D => n6344, Z => 
                           n6494);
   U6099 : NR2 port map( A => n6244, B => n6329, Z => n6344);
   U6100 : NR2 port map( A => n6291, B => n6329, Z => n6409);
   U6101 : ND2 port map( A => n4980, B => n6512, Z => n6511);
   U6102 : AO1 port map( A => n6426, B => n6281, C => n4982, D => n6513, Z => 
                           n6493);
   U6103 : AO6 port map( A => n6352, B => n6416, C => n4979, Z => n6513);
   U6104 : AO1 port map( A => n4994, B => n6514, C => n6515, D => n6516, Z => 
                           n6491);
   U6105 : AO4 port map( A => n6517, B => n4974, C => n6518, D => n6260, Z => 
                           n6516);
   U6106 : IV port map( A => n6519, Z => n6260);
   U6107 : AO1 port map( A => n6281, B => n6363, C => n6520, D => n6404, Z => 
                           n6518);
   U6108 : NR2 port map( A => n6363, B => n4979, Z => n6404);
   U6109 : AO4 port map( A => v_RAM_OUT0_26_port, B => n6244, C => n6329, D => 
                           n6427, Z => n6520);
   U6110 : IV port map( A => n6521, Z => n6363);
   U6111 : AO1 port map( A => n6408, B => n4359, C => n6522, D => n6523, Z => 
                           n6517);
   U6112 : AN3 port map( A => n6350, B => n6340, C => n6333, Z => n6523);
   U6113 : NR2 port map( A => v_RAM_OUT0_28_port, B => n6352, Z => n6522);
   U6114 : ND4 port map( A => n6524, B => n6525, C => n6526, D => n4971, Z => 
                           n6515);
   U6115 : ND4 port map( A => n6265, B => n6527, C => n6244, D => n4404, Z => 
                           n6526);
   U6116 : IV port map( A => n6276, Z => n6244);
   U6117 : ND3 port map( A => n6410, B => n6291, C => n6254, Z => n6525);
   U6118 : AO7 port map( A => n6528, B => n6292, C => n4978, Z => n6524);
   U6119 : NR3 port map( A => n4982, B => n4410, C => n6313, Z => n6528);
   U6120 : IV port map( A => n6529, Z => n6313);
   U6121 : AO3 port map( A => n6326, B => n6530, C => n6531, D => n6532, Z => 
                           n6514);
   U6122 : AO2 port map( A => n4975, B => n6533, C => n6534, D => n6265, Z => 
                           n6532);
   U6123 : ND2 port map( A => n6397, B => n6366, Z => n6533);
   U6124 : ND3 port map( A => n6267, B => n6382, C => n6333, Z => n6531);
   U6125 : ND2 port map( A => n6350, B => n6340, Z => n6530);
   U6126 : AO3 port map( A => n6535, B => n6444, C => n6536, D => n6537, Z => 
                           n4158);
   U6127 : AO6 port map( A => v_RAM_IN0_31_port, B => n6538, C => n6539, Z => 
                           n6537);
   U6128 : AO4 port map( A => n6540, B => n6541, C => n6542, D => n6543, Z => 
                           n6539);
   U6129 : EO port map( A => n6544, B => n6545, Z => n6542);
   U6130 : EN port map( A => n4931, B => n6546, Z => n6545);
   U6131 : EO port map( A => n6547, B => n6548, Z => n6540);
   U6132 : EO port map( A => n5821, B => n6549, Z => n6548);
   U6133 : AO2 port map( A => n6440, B => n6550, C => n6551, D => n6552, Z => 
                           n6536);
   U6134 : EN port map( A => n6553, B => n6554, Z => n6552);
   U6135 : EN port map( A => n4679, B => n6555, Z => n6554);
   U6136 : EO port map( A => v_KEY_COLUMN_31_port, B => v_DATA_COLUMN_31_port, 
                           Z => n6550);
   U6137 : EO port map( A => n6556, B => n6557, Z => n6535);
   U6138 : EN port map( A => n4775, B => n6558, Z => n6557);
   U6139 : MUX21H port map( A => t_STATE_RAM0_0_31_port, B => v_RAM_IN0_31_port
                           , S => n6480, Z => n4157);
   U6140 : MUX21H port map( A => t_STATE_RAM0_1_31_port, B => v_RAM_IN0_31_port
                           , S => n6481, Z => n4156);
   U6141 : MUX21H port map( A => t_STATE_RAM0_2_31_port, B => v_RAM_IN0_31_port
                           , S => n6482, Z => n4155);
   U6142 : MUX21H port map( A => t_STATE_RAM0_3_31_port, B => v_RAM_IN0_31_port
                           , S => n4498, Z => n4154);
   U6143 : AO3 port map( A => n6483, B => n4437, C => n6559, D => n6560, Z => 
                           n4153);
   U6144 : AO2 port map( A => t_STATE_RAM0_3_31_port, B => n6486, C => 
                           v_RAM_OUT0_31_port, D => n4513, Z => n6560);
   U6145 : AO2 port map( A => t_STATE_RAM0_1_31_port, B => n4564, C => 
                           t_STATE_RAM0_2_31_port, D => n4563, Z => n6559);
   U6146 : AO3 port map( A => n6437, B => n4372, C => n6561, D => n6562, Z => 
                           n4152);
   U6147 : AO6 port map( A => n6440, B => n6563, C => n6564, Z => n6562);
   U6148 : AO4 port map( A => n6565, B => n6444, C => n6566, D => n6446, Z => 
                           n6564);
   U6149 : EO port map( A => n6567, B => n6568, Z => n6566);
   U6150 : EN port map( A => n4707, B => n6553, Z => n6568);
   U6151 : EO port map( A => n6569, B => n6570, Z => n6553);
   U6152 : EO port map( A => n6571, B => n4712, Z => n6570);
   U6153 : EO port map( A => n6572, B => n6573, Z => n6565);
   U6154 : EN port map( A => n4834, B => n6558, Z => n6573);
   U6155 : EO port map( A => n6574, B => n6575, Z => n6558);
   U6156 : EO port map( A => n6576, B => n4838, Z => n6575);
   U6157 : EO port map( A => v_KEY_COLUMN_23_port, B => v_DATA_COLUMN_23_port, 
                           Z => n6563);
   U6158 : AO2 port map( A => n6462, B => n6577, C => n6464, D => n6578, Z => 
                           n6561);
   U6159 : EO port map( A => n6579, B => n6580, Z => n6578);
   U6160 : EN port map( A => n6229, B => n6549, Z => n6580);
   U6161 : EN port map( A => n6581, B => n6582, Z => n6549);
   U6162 : EN port map( A => n6583, B => n6584, Z => n6582);
   U6163 : EO port map( A => n6585, B => n6586, Z => n6577);
   U6164 : EN port map( A => n4950, B => n6544, Z => n6586);
   U6165 : EN port map( A => n6587, B => n6588, Z => n6544);
   U6166 : EO port map( A => n6589, B => n4954, Z => n6588);
   U6167 : MUX21L port map( A => n4421, B => n4372, S => n6480, Z => n4151);
   U6168 : MUX21H port map( A => t_STATE_RAM0_1_23_port, B => v_RAM_IN0_23_port
                           , S => n6481, Z => n4150);
   U6169 : MUX21H port map( A => t_STATE_RAM0_2_23_port, B => v_RAM_IN0_23_port
                           , S => n6482, Z => n4149);
   U6170 : MUX21H port map( A => t_STATE_RAM0_3_23_port, B => v_RAM_IN0_23_port
                           , S => n4498, Z => n4148);
   U6171 : AO3 port map( A => n6483, B => n4421, C => n6590, D => n6591, Z => 
                           n4147);
   U6172 : AO2 port map( A => t_STATE_RAM0_3_23_port, B => n6486, C => 
                           v_RAM_OUT0_23_port, D => n4513, Z => n6591);
   U6173 : AO2 port map( A => t_STATE_RAM0_1_23_port, B => n4564, C => 
                           t_STATE_RAM0_2_23_port, D => n4563, Z => n6590);
   U6174 : AO3 port map( A => n6592, B => n6444, C => n6593, D => n6594, Z => 
                           n4146);
   U6175 : AO6 port map( A => v_RAM_IN0_15_port, B => n6538, C => n6595, Z => 
                           n6594);
   U6176 : AO4 port map( A => n6596, B => n6541, C => n6597, D => n6543, Z => 
                           n6595);
   U6177 : EO port map( A => n6598, B => n6599, Z => n6597);
   U6178 : EO port map( A => n6600, B => n6601, Z => n6599);
   U6179 : EN port map( A => n4852, B => n6602, Z => n6598);
   U6180 : EO port map( A => n6603, B => n6604, Z => n6596);
   U6181 : EN port map( A => n6605, B => n6606, Z => n6604);
   U6182 : EN port map( A => n5008, B => n6607, Z => n6603);
   U6183 : AO2 port map( A => n6440, B => n6608, C => n6551, D => n6609, Z => 
                           n6593);
   U6184 : EO port map( A => n6610, B => n6611, Z => n6609);
   U6185 : EO port map( A => n6612, B => n6613, Z => n6611);
   U6186 : EN port map( A => n4583, B => n6614, Z => n6610);
   U6187 : EO port map( A => v_KEY_COLUMN_15_port, B => v_DATA_COLUMN_15_port, 
                           Z => n6608);
   U6188 : EO port map( A => n6615, B => n6616, Z => n6592);
   U6189 : EO port map( A => n6617, B => n6618, Z => n6616);
   U6190 : EN port map( A => n4734, B => n6619, Z => n6615);
   U6191 : MUX21H port map( A => t_STATE_RAM0_0_15_port, B => v_RAM_IN0_15_port
                           , S => n6480, Z => n4145);
   U6192 : MUX21H port map( A => t_STATE_RAM0_1_15_port, B => v_RAM_IN0_15_port
                           , S => n6481, Z => n4144);
   U6193 : MUX21H port map( A => t_STATE_RAM0_2_15_port, B => v_RAM_IN0_15_port
                           , S => n6482, Z => n4143);
   U6194 : MUX21H port map( A => t_STATE_RAM0_3_15_port, B => v_RAM_IN0_15_port
                           , S => n4498, Z => n4142);
   U6195 : AO3 port map( A => n6483, B => n4438, C => n6620, D => n6621, Z => 
                           n4141);
   U6196 : AO2 port map( A => t_STATE_RAM0_3_15_port, B => n6486, C => 
                           v_RAM_OUT0_15_port, D => n4513, Z => n6621);
   U6197 : AO2 port map( A => t_STATE_RAM0_1_15_port, B => n4564, C => 
                           t_STATE_RAM0_2_15_port, D => n4563, Z => n6620);
   U6198 : AO3 port map( A => n6622, B => n6444, C => n6623, D => n6624, Z => 
                           n4140);
   U6199 : AO6 port map( A => v_RAM_IN0_7_port, B => n6538, C => n6625, Z => 
                           n6624);
   U6200 : AO4 port map( A => n6626, B => n6541, C => n6627, D => n6543, Z => 
                           n6625);
   U6201 : EO port map( A => n6628, B => n6629, Z => n6627);
   U6202 : EN port map( A => n6630, B => n6601, Z => n6629);
   U6203 : EO port map( A => n6631, B => n6632, Z => n6601);
   U6204 : EN port map( A => n6589, B => n4918, Z => n6632);
   U6205 : EN port map( A => n6633, B => n6634, Z => n6589);
   U6206 : EN port map( A => n4857, B => n6635, Z => n6628);
   U6207 : EO port map( A => n6636, B => n6637, Z => n6626);
   U6208 : EN port map( A => n6638, B => n6606, Z => n6637);
   U6209 : EO port map( A => n6639, B => n6640, Z => n6606);
   U6210 : EO port map( A => n6583, B => n5507, Z => n6640);
   U6211 : EN port map( A => n6641, B => n6642, Z => n6583);
   U6212 : EN port map( A => n5095, B => n6643, Z => n6636);
   U6213 : AO2 port map( A => n6440, B => n6644, C => n6551, D => n6645, Z => 
                           n6623);
   U6214 : EO port map( A => n6646, B => n6647, Z => n6645);
   U6215 : EN port map( A => n6648, B => n6613, Z => n6647);
   U6216 : EN port map( A => n6649, B => n6650, Z => n6613);
   U6217 : EN port map( A => n6571, B => n4621, Z => n6650);
   U6218 : EN port map( A => n6651, B => n6652, Z => n6571);
   U6219 : EN port map( A => n4589, B => n6653, Z => n6646);
   U6220 : EO port map( A => v_KEY_COLUMN_7_port, B => v_DATA_COLUMN_7_port, Z 
                           => n6644);
   U6221 : EO port map( A => n6654, B => n6655, Z => n6622);
   U6222 : EN port map( A => n6656, B => n6618, Z => n6655);
   U6223 : EO port map( A => n6657, B => n6658, Z => n6618);
   U6224 : EN port map( A => n6576, B => n4760, Z => n6658);
   U6225 : EN port map( A => n6659, B => n6660, Z => n6576);
   U6226 : EN port map( A => n4739, B => n6661, Z => n6654);
   U6227 : MUX21H port map( A => t_STATE_RAM0_0_7_port, B => v_RAM_IN0_7_port, 
                           S => n6480, Z => n4139);
   U6228 : MUX21H port map( A => t_STATE_RAM0_1_7_port, B => v_RAM_IN0_7_port, 
                           S => n6481, Z => n4138);
   U6229 : MUX21H port map( A => t_STATE_RAM0_2_7_port, B => v_RAM_IN0_7_port, 
                           S => n6482, Z => n4137);
   U6230 : MUX21H port map( A => t_STATE_RAM0_3_7_port, B => v_RAM_IN0_7_port, 
                           S => n4498, Z => n4136);
   U6231 : AO3 port map( A => n6483, B => n4439, C => n6662, D => n6663, Z => 
                           n4135);
   U6232 : AO2 port map( A => t_STATE_RAM0_3_7_port, B => n6486, C => 
                           v_RAM_OUT0_7_port, D => n4513, Z => n6663);
   U6233 : AO2 port map( A => t_STATE_RAM0_1_7_port, B => n4564, C => 
                           t_STATE_RAM0_2_7_port, D => n4563, Z => n6662);
   U6234 : AO7 port map( A => n6664, B => n5009, C => n6665, Z => n4134);
   U6235 : AO2 port map( A => n6231, B => n4723, C => n7924, D => n6232, Z => 
                           n6665);
   U6236 : IV port map( A => n6666, Z => n4723);
   U6237 : AO7 port map( A => n6667, B => n6235, C => n6668, Z => n6666);
   U6238 : MUX21L port map( A => n6669, B => n6670, S => n4396, Z => n6668);
   U6239 : ND4 port map( A => n6671, B => n6672, C => n6673, D => n6674, Z => 
                           n6670);
   U6240 : AO2 port map( A => n4968, B => n6675, C => n6676, D => n6677, Z => 
                           n6674);
   U6241 : ND2 port map( A => n6427, B => n6416, Z => n6675);
   U6242 : IV port map( A => n6678, Z => n6673);
   U6243 : AO4 port map( A => n6679, B => n6350, C => n6362, D => n6680, Z => 
                           n6678);
   U6244 : EO1 port map( A => n6402, B => n6395, C => n4971, D => n6378, Z => 
                           n6672);
   U6245 : NR2 port map( A => n6381, B => n6290, Z => n6378);
   U6246 : ND2 port map( A => n6382, B => n6527, Z => n6395);
   U6247 : AO2 port map( A => n6254, B => n6681, C => n6292, D => n6264, Z => 
                           n6671);
   U6248 : NR4 port map( A => n6682, B => n6683, C => n6684, D => n6685, Z => 
                           n6669);
   U6249 : AO4 port map( A => n6686, B => n6687, C => n6240, D => n6370, Z => 
                           n6685);
   U6250 : AO3 port map( A => n6688, B => n6371, C => v_RAM_OUT0_29_port, D => 
                           n6689, Z => n6687);
   U6251 : EO1 port map( A => n6690, B => n6269, C => n6306, D => n6691, Z => 
                           n6689);
   U6252 : IV port map( A => n6249, Z => n6269);
   U6253 : NR2 port map( A => n4976, B => n6289, Z => n6249);
   U6254 : AO3 port map( A => n6692, B => n6300, C => n6693, D => n6694, Z => 
                           n6686);
   U6255 : AO2 port map( A => n6369, B => n6695, C => n6696, D => n6697, Z => 
                           n6694);
   U6256 : ND2 port map( A => n6410, B => n6506, Z => n6697);
   U6257 : ND2 port map( A => n4978, B => n6403, Z => n6695);
   U6258 : AO2 port map( A => n6698, B => n6359, C => n6699, D => n6700, Z => 
                           n6693);
   U6259 : NR2 port map( A => n4996, B => n6381, Z => n6698);
   U6260 : NR2 port map( A => n6701, B => n6277, Z => n6692);
   U6261 : AO4 port map( A => n6264, B => n6247, C => n6330, D => n6391, Z => 
                           n6684);
   U6262 : AO4 port map( A => n6270, B => n6278, C => n6680, D => n6702, Z => 
                           n6683);
   U6263 : AO3 port map( A => n6347, B => n6679, C => n6703, D => n6704, Z => 
                           n6682);
   U6264 : ND3 port map( A => n6397, B => n6366, C => n6677, Z => n6704);
   U6265 : OR3 port map( A => n6676, B => n6364, C => n4971, Z => n6703);
   U6266 : AO1 port map( A => n6705, B => n4978, C => n6706, D => n6707, Z => 
                           n6667);
   U6267 : AO4 port map( A => n6708, B => n6709, C => n6298, D => n6310, Z => 
                           n6707);
   U6268 : ND2 port map( A => n6506, B => n6263, Z => n6310);
   U6269 : AO6 port map( A => n6380, B => n6710, C => n6359, Z => n6708);
   U6270 : NR2 port map( A => n4364, B => v_RAM_OUT0_26_port, Z => n6380);
   U6271 : AO7 port map( A => n6309, B => n6291, C => n6711, Z => n6706);
   U6272 : AO2 port map( A => n6377, B => n6710, C => n6690, D => n6712, Z => 
                           n6711);
   U6273 : ND2 port map( A => n4980, B => n6350, Z => n6710);
   U6274 : AO7 port map( A => n6287, B => n6306, C => n6300, Z => n6705);
   U6275 : AO3 port map( A => n6437, B => n4373, C => n6713, D => n6714, Z => 
                           n4133);
   U6276 : AO6 port map( A => n6440, B => n6715, C => n6716, Z => n6714);
   U6277 : AO4 port map( A => n6717, B => n6444, C => n6718, D => n6446, Z => 
                           n6716);
   U6278 : EO port map( A => n6719, B => n6720, Z => n6718);
   U6279 : EN port map( A => n4715, B => n6721, Z => n6720);
   U6280 : EN port map( A => n4592, B => n4621, Z => n6719);
   U6281 : EO port map( A => n6722, B => n6723, Z => n6717);
   U6282 : EN port map( A => n4840, B => n6724, Z => n6723);
   U6283 : EN port map( A => n4741, B => n4760, Z => n6722);
   U6284 : EO port map( A => v_KEY_COLUMN_30_port, B => v_DATA_COLUMN_30_port, 
                           Z => n6715);
   U6285 : AO2 port map( A => n6462, B => n6725, C => n6464, D => n6726, Z => 
                           n6713);
   U6286 : EO port map( A => n6727, B => n6728, Z => n6726);
   U6287 : EN port map( A => n6383, B => n6729, Z => n6728);
   U6288 : EO port map( A => n5161, B => n5507, Z => n6727);
   U6289 : EO port map( A => n6730, B => n6731, Z => n6725);
   U6290 : EN port map( A => n4956, B => n6732, Z => n6731);
   U6291 : EN port map( A => n4859, B => n4918, Z => n6730);
   U6292 : MUX21L port map( A => n4422, B => n4373, S => n6480, Z => n4132);
   U6293 : MUX21H port map( A => t_STATE_RAM0_1_30_port, B => v_RAM_IN0_30_port
                           , S => n6481, Z => n4131);
   U6294 : MUX21H port map( A => t_STATE_RAM0_2_30_port, B => v_RAM_IN0_30_port
                           , S => n6482, Z => n4130);
   U6295 : MUX21H port map( A => t_STATE_RAM0_3_30_port, B => v_RAM_IN0_30_port
                           , S => n4498, Z => n4129);
   U6296 : AO3 port map( A => n6483, B => n4422, C => n6733, D => n6734, Z => 
                           n4128);
   U6297 : AO2 port map( A => t_STATE_RAM0_3_30_port, B => n6486, C => 
                           v_RAM_OUT0_30_port, D => n4513, Z => n6734);
   U6298 : AO2 port map( A => t_STATE_RAM0_1_30_port, B => n4564, C => 
                           t_STATE_RAM0_2_30_port, D => n4563, Z => n6733);
   U6299 : AO3 port map( A => n6437, B => n4374, C => n6735, D => n6736, Z => 
                           n4127);
   U6300 : AO6 port map( A => n6440, B => n6737, C => n6738, Z => n6736);
   U6301 : AO4 port map( A => n6739, B => n6444, C => n6740, D => n6446, Z => 
                           n6738);
   U6302 : EO port map( A => n6741, B => n6742, Z => n6740);
   U6303 : EN port map( A => n4715, B => n6743, Z => n6742);
   U6304 : EN port map( A => n4589, B => n4690, Z => n6741);
   U6305 : EO port map( A => n6744, B => n6745, Z => n6739);
   U6306 : EN port map( A => n4840, B => n6746, Z => n6745);
   U6307 : EN port map( A => n4739, B => n4783, Z => n6744);
   U6308 : EO port map( A => v_KEY_COLUMN_22_port, B => v_DATA_COLUMN_22_port, 
                           Z => n6737);
   U6309 : AO2 port map( A => n6462, B => n6747, C => n6464, D => n6748, Z => 
                           n6735);
   U6310 : EO port map( A => n6749, B => n6750, Z => n6748);
   U6311 : EN port map( A => n6383, B => n6751, Z => n6750);
   U6312 : EN port map( A => n5095, B => n6029, Z => n6749);
   U6313 : EO port map( A => n6752, B => n6753, Z => n6747);
   U6314 : EN port map( A => n4956, B => n6754, Z => n6753);
   U6315 : EN port map( A => n4857, B => n4939, Z => n6752);
   U6316 : MUX21L port map( A => n4423, B => n4374, S => n6480, Z => n4126);
   U6317 : MUX21H port map( A => t_STATE_RAM0_1_22_port, B => v_RAM_IN0_22_port
                           , S => n6481, Z => n4125);
   U6318 : MUX21H port map( A => t_STATE_RAM0_2_22_port, B => v_RAM_IN0_22_port
                           , S => n6482, Z => n4124);
   U6319 : MUX21H port map( A => t_STATE_RAM0_3_22_port, B => v_RAM_IN0_22_port
                           , S => n4498, Z => n4123);
   U6320 : AO3 port map( A => n6483, B => n4423, C => n6755, D => n6756, Z => 
                           n4122);
   U6321 : AO2 port map( A => t_STATE_RAM0_3_22_port, B => n6486, C => 
                           v_RAM_OUT0_22_port, D => n4513, Z => n6756);
   U6322 : AO2 port map( A => t_STATE_RAM0_1_22_port, B => n4564, C => 
                           t_STATE_RAM0_2_22_port, D => n4563, Z => n6755);
   U6323 : AO3 port map( A => n6437, B => n4375, C => n6757, D => n6758, Z => 
                           n4121);
   U6324 : AO6 port map( A => n6440, B => n6759, C => n6760, Z => n6758);
   U6325 : AO4 port map( A => n6761, B => n6444, C => n6762, D => n6446, Z => 
                           n6760);
   U6326 : EO port map( A => n6763, B => n6764, Z => n6762);
   U6327 : EN port map( A => n4712, B => n6721, Z => n6764);
   U6328 : EO port map( A => n6765, B => n6766, Z => n6721);
   U6329 : EN port map( A => n6767, B => n6651, Z => n6766);
   U6330 : EN port map( A => n4622, B => n4690, Z => n6763);
   U6331 : EO port map( A => n6768, B => n6769, Z => n6761);
   U6332 : EN port map( A => n4838, B => n6724, Z => n6769);
   U6333 : EO port map( A => n6770, B => n6771, Z => n6724);
   U6334 : EN port map( A => n6772, B => n6659, Z => n6771);
   U6335 : EN port map( A => n4761, B => n4783, Z => n6768);
   U6336 : EO port map( A => v_KEY_COLUMN_14_port, B => v_DATA_COLUMN_14_port, 
                           Z => n6759);
   U6337 : AO2 port map( A => n6462, B => n6773, C => n6464, D => n6774, Z => 
                           n6757);
   U6338 : EO port map( A => n6775, B => n6776, Z => n6774);
   U6339 : EN port map( A => n6315, B => n6729, Z => n6776);
   U6340 : EN port map( A => n6777, B => n6778, Z => n6729);
   U6341 : EN port map( A => n6779, B => n6641, Z => n6778);
   U6342 : EN port map( A => n5575, B => n6029, Z => n6775);
   U6343 : EO port map( A => n6780, B => n6781, Z => n6773);
   U6344 : EN port map( A => n4954, B => n6732, Z => n6781);
   U6345 : EN port map( A => n6782, B => n6783, Z => n6732);
   U6346 : EN port map( A => n6784, B => n6633, Z => n6783);
   U6347 : EN port map( A => n4919, B => n4939, Z => n6780);
   U6348 : MUX21L port map( A => n4424, B => n4375, S => n6480, Z => n4120);
   U6349 : MUX21H port map( A => t_STATE_RAM0_1_14_port, B => v_RAM_IN0_14_port
                           , S => n6481, Z => n4119);
   U6350 : MUX21H port map( A => t_STATE_RAM0_2_14_port, B => v_RAM_IN0_14_port
                           , S => n6482, Z => n4118);
   U6351 : MUX21H port map( A => t_STATE_RAM0_3_14_port, B => v_RAM_IN0_14_port
                           , S => n4498, Z => n4117);
   U6352 : AO3 port map( A => n6483, B => n4424, C => n6785, D => n6786, Z => 
                           n4116);
   U6353 : AO2 port map( A => t_STATE_RAM0_3_14_port, B => n6486, C => 
                           v_RAM_OUT0_14_port, D => n4513, Z => n6786);
   U6354 : AO2 port map( A => t_STATE_RAM0_1_14_port, B => n4564, C => 
                           t_STATE_RAM0_2_14_port, D => n4563, Z => n6785);
   U6355 : AO3 port map( A => n6437, B => n4376, C => n6787, D => n6788, Z => 
                           n4115);
   U6356 : AO6 port map( A => n6440, B => n6789, C => n6790, Z => n6788);
   U6357 : AO4 port map( A => n6791, B => n6444, C => n6792, D => n6446, Z => 
                           n6790);
   U6358 : EO port map( A => n6793, B => n6794, Z => n6792);
   U6359 : EN port map( A => n4684, B => n6743, Z => n6794);
   U6360 : EO port map( A => n6767, B => n6795, Z => n6743);
   U6361 : EN port map( A => n6449, B => n6796, Z => n6795);
   U6362 : EO port map( A => n6797, B => n6798, Z => n6767);
   U6363 : EN port map( A => n4592, B => n6799, Z => n6793);
   U6364 : EO port map( A => n6800, B => n6801, Z => n6791);
   U6365 : EN port map( A => n4779, B => n6746, Z => n6801);
   U6366 : EO port map( A => n6772, B => n6802, Z => n6746);
   U6367 : EN port map( A => n6461, B => n6803, Z => n6802);
   U6368 : EO port map( A => n6804, B => n6805, Z => n6772);
   U6369 : EN port map( A => n4741, B => n6806, Z => n6800);
   U6370 : EO port map( A => v_KEY_COLUMN_6_port, B => v_DATA_COLUMN_6_port, Z 
                           => n6789);
   U6371 : AO2 port map( A => n6462, B => n6807, C => n6464, D => n6808, Z => 
                           n6787);
   U6372 : EO port map( A => n6809, B => n6810, Z => n6808);
   U6373 : EN port map( A => n5907, B => n6751, Z => n6810);
   U6374 : EN port map( A => n6779, B => n6811, Z => n6751);
   U6375 : EN port map( A => n6812, B => n6813, Z => n6811);
   U6376 : EO port map( A => n6814, B => n6815, Z => n6779);
   U6377 : EN port map( A => n5161, B => n6816, Z => n6809);
   U6378 : EO port map( A => n6817, B => n6818, Z => n6807);
   U6379 : EN port map( A => n4935, B => n6754, Z => n6818);
   U6380 : EN port map( A => n6784, B => n6819, Z => n6754);
   U6381 : EN port map( A => n6477, B => n6820, Z => n6819);
   U6382 : EO port map( A => n6821, B => n6822, Z => n6784);
   U6383 : EN port map( A => n4859, B => n6823, Z => n6817);
   U6384 : MUX21L port map( A => n4425, B => n4376, S => n6480, Z => n4114);
   U6385 : MUX21H port map( A => t_STATE_RAM0_1_6_port, B => v_RAM_IN0_6_port, 
                           S => n6481, Z => n4113);
   U6386 : MUX21H port map( A => t_STATE_RAM0_2_6_port, B => v_RAM_IN0_6_port, 
                           S => n6482, Z => n4112);
   U6387 : MUX21H port map( A => t_STATE_RAM0_3_6_port, B => v_RAM_IN0_6_port, 
                           S => n4498, Z => n4111);
   U6388 : AO3 port map( A => n6483, B => n4425, C => n6824, D => n6825, Z => 
                           n4110);
   U6389 : AO2 port map( A => t_STATE_RAM0_3_6_port, B => n6486, C => 
                           v_RAM_OUT0_6_port, D => n4513, Z => n6825);
   U6390 : AO2 port map( A => t_STATE_RAM0_1_6_port, B => n4564, C => 
                           t_STATE_RAM0_2_6_port, D => n4563, Z => n6824);
   U6391 : AO7 port map( A => n6826, B => n5009, C => n6827, Z => n4109);
   U6392 : AO2 port map( A => n6231, B => n4726, C => n7930, D => n6232, Z => 
                           n6827);
   U6393 : MUX21L port map( A => n6828, B => n4966, S => n4396, Z => n4726);
   U6394 : ND4 port map( A => n6829, B => n6830, C => n6831, D => n6832, Z => 
                           n4966);
   U6395 : AO1 port map( A => n6519, B => n6833, C => n6834, D => n6835, Z => 
                           n6832);
   U6396 : AO4 port map( A => n6836, B => n6266, C => n6691, D => n4971, Z => 
                           n6835);
   U6397 : NR2 port map( A => n6837, B => n6277, Z => n6691);
   U6398 : IV port map( A => n4994, Z => n6266);
   U6399 : NR2 port map( A => n6838, B => n6839, Z => n6836);
   U6400 : AO4 port map( A => n6428, B => n6329, C => n6326, D => n6429, Z => 
                           n6839);
   U6401 : ND2 port map( A => n6688, B => n6416, Z => n6429);
   U6402 : EON1 port map( A => n6499, B => n4979, C => n6840, D => n6265, Z => 
                           n6838);
   U6403 : NR2 port map( A => n6289, B => n6676, Z => n6499);
   U6404 : AO4 port map( A => n6240, B => n6427, C => n6247, D => n6366, Z => 
                           n6834);
   U6405 : IV port map( A => n6841, Z => n6366);
   U6406 : IV port map( A => n4968, Z => n6247);
   U6407 : AO3 port map( A => n4979, B => n6505, C => n6433, D => n6842, Z => 
                           n6833);
   U6408 : AO2 port map( A => n6265, B => n6843, C => n6281, D => n6844, Z => 
                           n6842);
   U6409 : ND2 port map( A => n6416, B => n6413, Z => n6844);
   U6410 : ND2 port map( A => n6382, B => n6274, Z => n6843);
   U6411 : IV port map( A => n6336, Z => n6274);
   U6412 : AO2 port map( A => n6333, B => n6364, C => n6362, D => n4975, Z => 
                           n6433);
   U6413 : ND2 port map( A => n6505, B => n6275, Z => n6362);
   U6414 : AO2 port map( A => n6677, B => n6426, C => n6845, D => n6330, Z => 
                           n6831);
   U6415 : AO7 port map( A => n6402, B => n4968, C => n6846, Z => n6830);
   U6416 : AO2 port map( A => n6847, B => n6254, C => n6253, D => n6848, Z => 
                           n6829);
   U6417 : ND2 port map( A => n6240, B => n6680, Z => n6848);
   U6418 : NR2 port map( A => n6367, B => n6529, Z => n6847);
   U6419 : AO3 port map( A => n6849, B => n4971, C => n6850, D => n6851, Z => 
                           n6828);
   U6420 : AO2 port map( A => n6252, B => n4983, C => v_RAM_OUT0_29_port, D => 
                           n4981, Z => n6851);
   U6421 : ND4 port map( A => n6852, B => n6853, C => n6854, D => n6855, Z => 
                           n4981);
   U6422 : AO2 port map( A => n6856, B => n6690, C => n6696, D => n6857, Z => 
                           n6855);
   U6423 : ND2 port map( A => n6293, B => n6413, Z => n6857);
   U6424 : IV port map( A => n6676, Z => n6413);
   U6425 : NR2 port map( A => n4368, B => v_RAM_OUT0_24_port, Z => n6676);
   U6426 : NR2 port map( A => n6841, B => n4967, Z => n6856);
   U6427 : AO2 port map( A => n6365, B => n6858, C => n6700, D => n6323, Z => 
                           n6854);
   U6428 : ND2 port map( A => n6350, B => n6339, Z => n6323);
   U6429 : AO2 port map( A => n6359, B => n6293, C => n6368, D => n6427, Z => 
                           n6853);
   U6430 : AO2 port map( A => n6377, B => n6264, C => n6369, D => n6370, Z => 
                           n6852);
   U6431 : AO3 port map( A => n5004, B => n4978, C => n6859, D => n6860, Z => 
                           n4983);
   U6432 : AO2 port map( A => n6336, B => n6333, C => n6861, D => n4975, Z => 
                           n6860);
   U6433 : NR2 port map( A => n6403, B => v_RAM_OUT0_24_port, Z => n6336);
   U6434 : ND2 port map( A => n6265, B => n6352, Z => n6859);
   U6435 : AO2 port map( A => n4968, B => n6862, C => n6250, D => n6863, Z => 
                           n6850);
   U6436 : AO3 port map( A => n6329, B => n4976, C => n6864, D => n6434, Z => 
                           n6863);
   U6437 : IV port map( A => n6348, Z => n6434);
   U6438 : NR2 port map( A => n6506, B => n4979, Z => n6348);
   U6439 : ND2 port map( A => n6346, B => n6333, Z => n6864);
   U6440 : ND2 port map( A => n6263, B => n6527, Z => n6862);
   U6441 : IV port map( A => n6299, Z => n6527);
   U6442 : IV port map( A => n6346, Z => n6263);
   U6443 : AO3 port map( A => n6865, B => n6444, C => n6866, D => n6867, Z => 
                           n4108);
   U6444 : AO6 port map( A => v_RAM_IN0_21_port, B => n6538, C => n6868, Z => 
                           n6867);
   U6445 : AO4 port map( A => n6869, B => n6541, C => n6870, D => n6543, Z => 
                           n6868);
   U6446 : EO port map( A => n6871, B => n6872, Z => n6870);
   U6447 : EN port map( A => n6873, B => n6874, Z => n6872);
   U6448 : EN port map( A => n4958, B => n6875, Z => n6871);
   U6449 : EO port map( A => n4859, B => n4940, Z => n6875);
   U6450 : EO port map( A => n6876, B => n6877, Z => n6869);
   U6451 : EN port map( A => n6878, B => n6879, Z => n6877);
   U6452 : EO port map( A => n6490, B => n6880, Z => n6876);
   U6453 : EO port map( A => n5161, B => n6030, Z => n6880);
   U6454 : AO2 port map( A => n6440, B => n6881, C => n6551, D => n6882, Z => 
                           n6866);
   U6455 : EO port map( A => n6883, B => n6884, Z => n6882);
   U6456 : EN port map( A => n6885, B => n6886, Z => n6884);
   U6457 : EN port map( A => n4718, B => n6887, Z => n6883);
   U6458 : EO port map( A => n4592, B => n4691, Z => n6887);
   U6459 : EO port map( A => v_KEY_COLUMN_21_port, B => v_DATA_COLUMN_21_port, 
                           Z => n6881);
   U6460 : EO port map( A => n6888, B => n6889, Z => n6865);
   U6461 : EN port map( A => n6890, B => n6891, Z => n6889);
   U6462 : EN port map( A => n4842, B => n6892, Z => n6888);
   U6463 : EO port map( A => n4741, B => n4784, Z => n6892);
   U6464 : MUX21H port map( A => t_STATE_RAM0_0_21_port, B => v_RAM_IN0_21_port
                           , S => n6480, Z => n4107);
   U6465 : MUX21H port map( A => t_STATE_RAM0_1_21_port, B => v_RAM_IN0_21_port
                           , S => n6481, Z => n4106);
   U6466 : MUX21H port map( A => t_STATE_RAM0_2_21_port, B => v_RAM_IN0_21_port
                           , S => n6482, Z => n4105);
   U6467 : MUX21H port map( A => t_STATE_RAM0_3_21_port, B => v_RAM_IN0_21_port
                           , S => n4498, Z => n4104);
   U6468 : AO3 port map( A => n6483, B => n4440, C => n6893, D => n6894, Z => 
                           n4103);
   U6469 : AO2 port map( A => t_STATE_RAM0_3_21_port, B => n6486, C => 
                           v_RAM_OUT0_21_port, D => n4513, Z => n6894);
   U6470 : AO2 port map( A => t_STATE_RAM0_1_21_port, B => n4564, C => 
                           t_STATE_RAM0_2_21_port, D => n4563, Z => n6893);
   U6471 : AO3 port map( A => n6895, B => n6444, C => n6896, D => n6897, Z => 
                           n4102);
   U6472 : AO6 port map( A => v_RAM_IN0_13_port, B => n6538, C => n6898, Z => 
                           n6897);
   U6473 : AO4 port map( A => n6899, B => n6541, C => n6900, D => n6543, Z => 
                           n6898);
   U6474 : EO port map( A => n6901, B => n6902, Z => n6900);
   U6475 : EN port map( A => n6874, B => n6903, Z => n6902);
   U6476 : EN port map( A => n4956, B => n6904, Z => n6901);
   U6477 : EO port map( A => n4921, B => n4940, Z => n6904);
   U6478 : EO port map( A => n6905, B => n6906, Z => n6899);
   U6479 : EN port map( A => n6878, B => n6907, Z => n6906);
   U6480 : EN port map( A => n6383, B => n6908, Z => n6905);
   U6481 : EO port map( A => n5624, B => n6030, Z => n6908);
   U6482 : AO2 port map( A => n6440, B => n6909, C => n6551, D => n6910, Z => 
                           n6896);
   U6483 : EO port map( A => n6911, B => n6912, Z => n6910);
   U6484 : EN port map( A => n6886, B => n6913, Z => n6912);
   U6485 : EN port map( A => n4715, B => n6914, Z => n6911);
   U6486 : EO port map( A => n4625, B => n4691, Z => n6914);
   U6487 : EO port map( A => v_KEY_COLUMN_13_port, B => v_DATA_COLUMN_13_port, 
                           Z => n6909);
   U6488 : EO port map( A => n6915, B => n6916, Z => n6895);
   U6489 : EN port map( A => n6891, B => n6917, Z => n6916);
   U6490 : EN port map( A => n4840, B => n6918, Z => n6915);
   U6491 : EO port map( A => n4763, B => n4784, Z => n6918);
   U6492 : MUX21H port map( A => t_STATE_RAM0_0_13_port, B => v_RAM_IN0_13_port
                           , S => n6480, Z => n4101);
   U6493 : MUX21H port map( A => t_STATE_RAM0_1_13_port, B => v_RAM_IN0_13_port
                           , S => n6481, Z => n4100);
   U6494 : MUX21H port map( A => t_STATE_RAM0_2_13_port, B => v_RAM_IN0_13_port
                           , S => n6482, Z => n4099);
   U6495 : MUX21H port map( A => t_STATE_RAM0_3_13_port, B => v_RAM_IN0_13_port
                           , S => n4498, Z => n4098);
   U6496 : AO3 port map( A => n6483, B => n4441, C => n6919, D => n6920, Z => 
                           n4097);
   U6497 : AO2 port map( A => t_STATE_RAM0_3_13_port, B => n6486, C => 
                           v_RAM_OUT0_13_port, D => n4513, Z => n6920);
   U6498 : AO2 port map( A => t_STATE_RAM0_1_13_port, B => n4564, C => 
                           t_STATE_RAM0_2_13_port, D => n4563, Z => n6919);
   U6499 : AO3 port map( A => n6921, B => n6444, C => n6922, D => n6923, Z => 
                           n4096);
   U6500 : AO6 port map( A => v_RAM_IN0_29_port, B => n6538, C => n6924, Z => 
                           n6923);
   U6501 : AO4 port map( A => n6925, B => n6541, C => n6926, D => n6543, Z => 
                           n6924);
   U6502 : EO port map( A => n6927, B => n6928, Z => n6926);
   U6503 : EO port map( A => n6903, B => n6929, Z => n6928);
   U6504 : EO port map( A => n6822, B => n6930, Z => n6903);
   U6505 : EO port map( A => n6931, B => n6932, Z => n6822);
   U6506 : EN port map( A => n4919, B => n6933, Z => n6927);
   U6507 : EO port map( A => n6934, B => n6935, Z => n6925);
   U6508 : EO port map( A => n6907, B => n6936, Z => n6935);
   U6509 : EO port map( A => n6815, B => n6937, Z => n6907);
   U6510 : EO port map( A => n6938, B => n6939, Z => n6815);
   U6511 : EN port map( A => n5575, B => n6490, Z => n6934);
   U6512 : AO2 port map( A => n6440, B => n6940, C => n6551, D => n6941, Z => 
                           n6922);
   U6513 : EO port map( A => n6942, B => n6943, Z => n6941);
   U6514 : EO port map( A => n6913, B => n6944, Z => n6943);
   U6515 : EN port map( A => n6798, B => n6648, Z => n6913);
   U6516 : EO port map( A => n6945, B => n6946, Z => n6798);
   U6517 : EN port map( A => n4622, B => n6947, Z => n6942);
   U6518 : EO port map( A => v_KEY_COLUMN_29_port, B => v_DATA_COLUMN_29_port, 
                           Z => n6940);
   U6519 : EO port map( A => n6948, B => n6949, Z => n6921);
   U6520 : EO port map( A => n6917, B => n6950, Z => n6949);
   U6521 : EO port map( A => n6805, B => n6951, Z => n6917);
   U6522 : EO port map( A => n6952, B => n6953, Z => n6805);
   U6523 : EN port map( A => n4761, B => n6954, Z => n6948);
   U6524 : MUX21H port map( A => t_STATE_RAM0_0_29_port, B => v_RAM_IN0_29_port
                           , S => n6480, Z => n4095);
   U6525 : MUX21H port map( A => t_STATE_RAM0_1_29_port, B => v_RAM_IN0_29_port
                           , S => n6481, Z => n4094);
   U6526 : MUX21H port map( A => t_STATE_RAM0_2_29_port, B => v_RAM_IN0_29_port
                           , S => n6482, Z => n4093);
   U6527 : MUX21H port map( A => t_STATE_RAM0_3_29_port, B => v_RAM_IN0_29_port
                           , S => n4498, Z => n4092);
   U6528 : AO3 port map( A => n6483, B => n4442, C => n6955, D => n6956, Z => 
                           n4091);
   U6529 : AO2 port map( A => t_STATE_RAM0_3_29_port, B => n6486, C => 
                           v_RAM_OUT0_29_port, D => n4513, Z => n6956);
   U6530 : AO2 port map( A => t_STATE_RAM0_1_29_port, B => n4564, C => 
                           t_STATE_RAM0_2_29_port, D => n4563, Z => n6955);
   U6531 : AO3 port map( A => n6957, B => n6444, C => n6958, D => n6959, Z => 
                           n4090);
   U6532 : AO6 port map( A => v_RAM_IN0_5_port, B => n6538, C => n6960, Z => 
                           n6959);
   U6533 : AO4 port map( A => n6961, B => n6541, C => n6962, D => n6543, Z => 
                           n6960);
   U6534 : EO port map( A => n6963, B => n6964, Z => n6962);
   U6535 : EO port map( A => n6873, B => n6929, Z => n6964);
   U6536 : EN port map( A => n6965, B => n6874, Z => n6929);
   U6537 : EO port map( A => n6966, B => n6967, Z => n6874);
   U6538 : IV port map( A => n6968, Z => n6966);
   U6539 : EO port map( A => n6821, B => n6600, Z => n6873);
   U6540 : EO port map( A => n6969, B => n6970, Z => n6821);
   U6541 : EN port map( A => n4921, B => n4939, Z => n6963);
   U6542 : EO port map( A => n6971, B => n6972, Z => n6961);
   U6543 : EO port map( A => n6879, B => n6936, Z => n6972);
   U6544 : EN port map( A => n6973, B => n6878, Z => n6936);
   U6545 : EO port map( A => n6974, B => n6975, Z => n6878);
   U6546 : IV port map( A => n6976, Z => n6974);
   U6547 : EO port map( A => n6814, B => n6977, Z => n6879);
   U6548 : EO port map( A => n6978, B => n6979, Z => n6814);
   U6549 : EN port map( A => n5624, B => n6029, Z => n6971);
   U6550 : AO2 port map( A => n6440, B => n6980, C => n6551, D => n6981, Z => 
                           n6958);
   U6551 : EO port map( A => n6982, B => n6983, Z => n6981);
   U6552 : EO port map( A => n6885, B => n6944, Z => n6983);
   U6553 : EN port map( A => n6984, B => n6886, Z => n6944);
   U6554 : EN port map( A => n6985, B => n6986, Z => n6886);
   U6555 : EO port map( A => n6797, B => n6612, Z => n6885);
   U6556 : EO port map( A => n6987, B => n6988, Z => n6797);
   U6557 : EN port map( A => n4625, B => n4690, Z => n6982);
   U6558 : EO port map( A => v_KEY_COLUMN_5_port, B => v_DATA_COLUMN_5_port, Z 
                           => n6980);
   U6559 : EO port map( A => n6989, B => n6990, Z => n6957);
   U6560 : EO port map( A => n6890, B => n6950, Z => n6990);
   U6561 : EN port map( A => n6991, B => n6891, Z => n6950);
   U6562 : EO port map( A => n6992, B => n6993, Z => n6891);
   U6563 : IV port map( A => n6994, Z => n6992);
   U6564 : EO port map( A => n6804, B => n6617, Z => n6890);
   U6565 : EO port map( A => n6995, B => n6996, Z => n6804);
   U6566 : EN port map( A => n4763, B => n4783, Z => n6989);
   U6567 : MUX21H port map( A => t_STATE_RAM0_0_5_port, B => v_RAM_IN0_5_port, 
                           S => n6480, Z => n4089);
   U6568 : MUX21H port map( A => t_STATE_RAM0_1_5_port, B => v_RAM_IN0_5_port, 
                           S => n6481, Z => n4088);
   U6569 : MUX21H port map( A => t_STATE_RAM0_2_5_port, B => v_RAM_IN0_5_port, 
                           S => n6482, Z => n4087);
   U6570 : MUX21H port map( A => t_STATE_RAM0_3_5_port, B => v_RAM_IN0_5_port, 
                           S => n4498, Z => n4086);
   U6571 : AO3 port map( A => n6483, B => n4443, C => n6997, D => n6998, Z => 
                           n4085);
   U6572 : AO2 port map( A => t_STATE_RAM0_3_5_port, B => n6486, C => 
                           v_RAM_OUT0_5_port, D => n4513, Z => n6998);
   U6573 : AO2 port map( A => t_STATE_RAM0_1_5_port, B => n4564, C => 
                           t_STATE_RAM0_2_5_port, D => n4563, Z => n6997);
   U6574 : AO3 port map( A => n6999, B => n6444, C => n7000, D => n7001, Z => 
                           n4084);
   U6575 : AO6 port map( A => v_RAM_IN0_2_port, B => n6538, C => n7002, Z => 
                           n7001);
   U6576 : AO4 port map( A => n7003, B => n6541, C => n7004, D => n6543, Z => 
                           n7002);
   U6577 : EO port map( A => n7005, B => n7006, Z => n7004);
   U6578 : EN port map( A => n7007, B => n7008, Z => n7006);
   U6579 : EN port map( A => n4927, B => n7009, Z => n7005);
   U6580 : EO port map( A => n4888, B => n4925, Z => n7009);
   U6581 : EO port map( A => n7010, B => n7011, Z => n7003);
   U6582 : EN port map( A => n7012, B => n7013, Z => n7011);
   U6583 : EN port map( A => n5756, B => n7014, Z => n7010);
   U6584 : EO port map( A => n5345, B => n5713, Z => n7014);
   U6585 : AO2 port map( A => n6440, B => n7015, C => n6551, D => n7016, Z => 
                           n7000);
   U6586 : EO port map( A => n7017, B => n7018, Z => n7016);
   U6587 : EO port map( A => n7019, B => n7020, Z => n7018);
   U6588 : EN port map( A => n4652, B => n7021, Z => n7017);
   U6589 : EO port map( A => n4604, B => n4631, Z => n7021);
   U6590 : EO port map( A => v_KEY_COLUMN_2_port, B => v_DATA_COLUMN_2_port, Z 
                           => n7015);
   U6591 : EO port map( A => n7022, B => n7023, Z => n6999);
   U6592 : EN port map( A => n7024, B => n7025, Z => n7023);
   U6593 : EN port map( A => n4770, B => n7026, Z => n7022);
   U6594 : EO port map( A => n4749, B => n4767, Z => n7026);
   U6595 : MUX21H port map( A => t_STATE_RAM0_0_2_port, B => v_RAM_IN0_2_port, 
                           S => n6480, Z => n4083);
   U6596 : MUX21H port map( A => t_STATE_RAM0_1_2_port, B => v_RAM_IN0_2_port, 
                           S => n6481, Z => n4082);
   U6597 : MUX21H port map( A => t_STATE_RAM0_2_2_port, B => v_RAM_IN0_2_port, 
                           S => n6482, Z => n4081);
   U6598 : MUX21H port map( A => t_STATE_RAM0_3_2_port, B => v_RAM_IN0_2_port, 
                           S => n4498, Z => n4080);
   U6599 : AO3 port map( A => n6483, B => n4444, C => n7027, D => n7028, Z => 
                           n4079);
   U6600 : AO2 port map( A => t_STATE_RAM0_3_2_port, B => n6486, C => 
                           v_RAM_OUT0_2_port, D => n4513, Z => n7028);
   U6601 : AO2 port map( A => t_STATE_RAM0_1_2_port, B => n4564, C => 
                           t_STATE_RAM0_2_2_port, D => n4563, Z => n7027);
   U6602 : AO7 port map( A => n7029, B => n5009, C => n7030, Z => n4078);
   U6603 : AO2 port map( A => n6231, B => n4729, C => n7936, D => n6232, Z => 
                           n7030);
   U6604 : IV port map( A => n7031, Z => n4729);
   U6605 : AO7 port map( A => n7032, B => n6235, C => n7033, Z => n7031);
   U6606 : MUX21L port map( A => n7034, B => n7035, S => n4396, Z => n7033);
   U6607 : ND4 port map( A => n7036, B => n7037, C => n7038, D => n7039, Z => 
                           n7035);
   U6608 : AO2 port map( A => n6699, B => n6845, C => n6402, D => n7040, Z => 
                           n7039);
   U6609 : ND2 port map( A => n6688, B => n6341, Z => n7040);
   U6610 : NR2 port map( A => n6347, B => n6837, Z => n6699);
   U6611 : AO2 port map( A => n6254, B => n7041, C => n6677, D => n6398, Z => 
                           n7038);
   U6612 : NR2 port map( A => n4974, B => n4979, Z => n6677);
   U6613 : ND2 port map( A => n6410, B => n6264, Z => n7041);
   U6614 : IV port map( A => n6277, Z => n6264);
   U6615 : EO1 port map( A => n6243, B => n6702, C => n6240, D => n6271, Z => 
                           n7037);
   U6616 : NR2 port map( A => n6277, B => n6841, Z => n6271);
   U6617 : ND2 port map( A => n6427, B => n6512, Z => n6702);
   U6618 : IV port map( A => n6701, Z => n6512);
   U6619 : AO2 port map( A => n7042, B => n6427, C => n4968, D => n6681, Z => 
                           n7036);
   U6620 : IV port map( A => n6303, Z => n6681);
   U6621 : NR4 port map( A => n7043, B => n7044, C => n7045, D => n7046, Z => 
                           n7034);
   U6622 : AO4 port map( A => n7047, B => n7048, C => n6240, D => n6408, Z => 
                           n7046);
   U6623 : OR2 port map( A => n6426, B => n6841, Z => n6408);
   U6624 : AO3 port map( A => n6306, B => n7049, C => v_RAM_OUT0_29_port, D => 
                           n7050, Z => n7048);
   U6625 : AO2 port map( A => n6369, B => n4972, C => n6368, D => n6352, Z => 
                           n7050);
   U6626 : IV port map( A => n6849, Z => n4972);
   U6627 : NR2 port map( A => n4976, B => n6364, Z => n6849);
   U6628 : AO3 port map( A => n6302, B => n6341, C => n7051, D => n7052, Z => 
                           n7047);
   U6629 : EO1 port map( A => n6690, B => v_RAM_OUT0_27_port, C => n6291, D => 
                           n6311, Z => n7052);
   U6630 : EO1 port map( A => n7053, B => n6696, C => n6371, D => n6305, Z => 
                           n7051);
   U6631 : NR2 port map( A => n6426, B => n6276, Z => n6305);
   U6632 : IV port map( A => n6377, Z => n6371);
   U6633 : NR2 port map( A => n6330, B => n6837, Z => n7053);
   U6634 : MUX21L port map( A => n6679, B => n7054, S => n6278, Z => n7045);
   U6635 : NR2 port map( A => n7055, B => n4968, Z => n7054);
   U6636 : NR2 port map( A => n4974, B => n6326, Z => n4968);
   U6637 : AN3 port map( A => n4967, B => v_RAM_OUT0_26_port, C => n6250, Z => 
                           n7055);
   U6638 : IV port map( A => n6845, Z => n6679);
   U6639 : NR2 port map( A => n4982, B => n4979, Z => n6845);
   U6640 : AO4 port map( A => n6391, B => n6251, C => n6534, D => n6270, Z => 
                           n7044);
   U6641 : IV port map( A => n6402, Z => n6270);
   U6642 : NR2 port map( A => n4982, B => n6337, Z => n6402);
   U6643 : NR2 port map( A => n6287, B => n6841, Z => n6534);
   U6644 : NR2 port map( A => n4976, B => n4355, Z => n6841);
   U6645 : ND2 port map( A => n6314, B => n6397, Z => n6251);
   U6646 : IV port map( A => n6254, Z => n6391);
   U6647 : AO4 port map( A => n6680, B => n4980, C => n4971, D => n7056, Z => 
                           n7043);
   U6648 : ND2 port map( A => n6382, B => n6267, Z => n7056);
   U6649 : IV port map( A => n6861, Z => n6267);
   U6650 : IV port map( A => n6253, Z => n6382);
   U6651 : IV port map( A => n7042, Z => n4971);
   U6652 : NR2 port map( A => n4974, B => n6337, Z => n7042);
   U6653 : IV port map( A => n6243, Z => n6680);
   U6654 : NR2 port map( A => n4974, B => n6329, Z => n6243);
   U6655 : IV port map( A => n6250, Z => n4974);
   U6656 : ND2 port map( A => v_RAM_OUT0_29_port, B => n4396, Z => n6235);
   U6657 : NR4 port map( A => n7057, B => n7058, C => n7059, D => n7060, Z => 
                           n7032);
   U6658 : AO4 port map( A => n6304, B => n6507, C => n6303, D => n6302, Z => 
                           n7060);
   U6659 : IV port map( A => n6359, Z => n6302);
   U6660 : NR2 port map( A => n6701, B => n6529, Z => n6303);
   U6661 : NR2 port map( A => v_RAM_OUT0_24_port, B => n6288, Z => n6529);
   U6662 : IV port map( A => n5005, Z => n6507);
   U6663 : IV port map( A => n6690, Z => n6304);
   U6664 : EON1 port map( A => n6298, B => n6858, C => n6284, D => n6377, Z => 
                           n7059);
   U6665 : IV port map( A => n6369, Z => n6298);
   U6666 : EON1 port map( A => n7061, B => n6306, C => n6414, D => n6700, Z => 
                           n7058);
   U6667 : ND2 port map( A => n6397, B => n6275, Z => n6414);
   U6668 : IV port map( A => n4967, Z => n6397);
   U6669 : IV port map( A => n6365, Z => n6306);
   U6670 : NR2 port map( A => n6277, B => n4996, Z => n7061);
   U6671 : AO4 port map( A => n7062, B => n6300, C => n6309, D => n7063, Z => 
                           n7057);
   U6672 : ND2 port map( A => n6416, B => n6352, Z => n7063);
   U6673 : IV port map( A => n6364, Z => n6416);
   U6674 : NR2 port map( A => n4355, B => n6288, Z => n6364);
   U6675 : IV port map( A => n6696, Z => n6309);
   U6676 : NR2 port map( A => n6861, B => n6239, Z => n7062);
   U6677 : NR2 port map( A => n6688, B => v_RAM_OUT0_24_port, Z => n6861);
   U6678 : AO3 port map( A => n7064, B => n6444, C => n7065, D => n7066, Z => 
                           n4077);
   U6679 : AO6 port map( A => v_RAM_IN0_18_port, B => n6538, C => n7067, Z => 
                           n7066);
   U6680 : AO4 port map( A => n7068, B => n6541, C => n7069, D => n6543, Z => 
                           n7067);
   U6681 : EO port map( A => n7070, B => n7071, Z => n7069);
   U6682 : EN port map( A => n7007, B => n7072, Z => n7071);
   U6683 : EO port map( A => n7073, B => n6479, Z => n7007);
   U6684 : EN port map( A => n4984, B => n7074, Z => n7070);
   U6685 : EN port map( A => n4946, B => n7075, Z => n7074);
   U6686 : EO port map( A => n7076, B => n7077, Z => n7068);
   U6687 : EO port map( A => n7029, B => n7078, Z => n7077);
   U6688 : EO port map( A => n7012, B => n7079, Z => n7076);
   U6689 : EN port map( A => n6164, B => n7080, Z => n7079);
   U6690 : EO port map( A => n7081, B => n7082, Z => n7012);
   U6691 : AO2 port map( A => n6440, B => n7083, C => n6551, D => n7084, Z => 
                           n7065);
   U6692 : EO port map( A => n7085, B => n7086, Z => n7084);
   U6693 : EO port map( A => n7019, B => n7087, Z => n7086);
   U6694 : EO port map( A => n7088, B => n6453, Z => n7019);
   U6695 : EN port map( A => n4727, B => n7089, Z => n7085);
   U6696 : EN port map( A => n4700, B => n7090, Z => n7089);
   U6697 : EO port map( A => v_KEY_COLUMN_18_port, B => v_DATA_COLUMN_18_port, 
                           Z => n7083);
   U6698 : EO port map( A => n7091, B => n7092, Z => n7064);
   U6699 : EN port map( A => n7024, B => n7093, Z => n7092);
   U6700 : EO port map( A => n7094, B => n6456, Z => n7024);
   U6701 : EN port map( A => n4848, B => n7095, Z => n7091);
   U6702 : EN port map( A => n4810, B => n7096, Z => n7095);
   U6703 : MUX21H port map( A => t_STATE_RAM0_0_18_port, B => v_RAM_IN0_18_port
                           , S => n6480, Z => n4076);
   U6704 : MUX21H port map( A => t_STATE_RAM0_1_18_port, B => v_RAM_IN0_18_port
                           , S => n6481, Z => n4075);
   U6705 : MUX21H port map( A => t_STATE_RAM0_2_18_port, B => v_RAM_IN0_18_port
                           , S => n6482, Z => n4074);
   U6706 : MUX21H port map( A => t_STATE_RAM0_3_18_port, B => v_RAM_IN0_18_port
                           , S => n4498, Z => n4073);
   U6707 : AO3 port map( A => n6483, B => n4445, C => n7097, D => n7098, Z => 
                           n4072);
   U6708 : AO2 port map( A => t_STATE_RAM0_3_18_port, B => n6486, C => 
                           v_RAM_OUT0_18_port, D => n4513, Z => n7098);
   U6709 : AO2 port map( A => t_STATE_RAM0_1_18_port, B => n4564, C => 
                           t_STATE_RAM0_2_18_port, D => n4563, Z => n7097);
   U6710 : AO3 port map( A => n7099, B => n6444, C => n7100, D => n7101, Z => 
                           n4071);
   U6711 : AO6 port map( A => v_RAM_IN0_9_port, B => n6538, C => n7102, Z => 
                           n7101);
   U6712 : AO4 port map( A => n7103, B => n6541, C => n7104, D => n6543, Z => 
                           n7102);
   U6713 : EO port map( A => n7105, B => n7106, Z => n7104);
   U6714 : EN port map( A => n7107, B => n7108, Z => n7106);
   U6715 : EN port map( A => n4946, B => n7109, Z => n7105);
   U6716 : EO port map( A => n7110, B => n7111, Z => n7103);
   U6717 : EN port map( A => n7112, B => n7113, Z => n7111);
   U6718 : EN port map( A => n6164, B => n7114, Z => n7110);
   U6719 : AO2 port map( A => n6440, B => n7115, C => n6551, D => n7116, Z => 
                           n7100);
   U6720 : EO port map( A => n7117, B => n7118, Z => n7116);
   U6721 : EO port map( A => n7119, B => n7120, Z => n7118);
   U6722 : EN port map( A => n4700, B => n7121, Z => n7117);
   U6723 : EO port map( A => v_KEY_COLUMN_9_port, B => v_DATA_COLUMN_9_port, Z 
                           => n7115);
   U6724 : EO port map( A => n7122, B => n7123, Z => n7099);
   U6725 : EN port map( A => n7124, B => n7125, Z => n7123);
   U6726 : EN port map( A => n4810, B => n7126, Z => n7122);
   U6727 : MUX21H port map( A => t_STATE_RAM0_0_9_port, B => v_RAM_IN0_9_port, 
                           S => n6480, Z => n4070);
   U6728 : MUX21H port map( A => t_STATE_RAM0_1_9_port, B => v_RAM_IN0_9_port, 
                           S => n6481, Z => n4069);
   U6729 : MUX21H port map( A => t_STATE_RAM0_2_9_port, B => v_RAM_IN0_9_port, 
                           S => n6482, Z => n4068);
   U6730 : MUX21H port map( A => t_STATE_RAM0_3_9_port, B => v_RAM_IN0_9_port, 
                           S => n4498, Z => n4067);
   U6731 : AO3 port map( A => n6483, B => n4446, C => n7127, D => n7128, Z => 
                           n4066);
   U6732 : AO2 port map( A => t_STATE_RAM0_3_9_port, B => n6486, C => 
                           v_RAM_OUT0_9_port, D => n4513, Z => n7128);
   U6733 : AO2 port map( A => t_STATE_RAM0_1_9_port, B => n4564, C => 
                           t_STATE_RAM0_2_9_port, D => n4563, Z => n7127);
   U6734 : AO3 port map( A => n7129, B => n6444, C => n7130, D => n7131, Z => 
                           n4065);
   U6735 : AO6 port map( A => v_RAM_IN0_28_port, B => n6538, C => n7132, Z => 
                           n7131);
   U6736 : AO4 port map( A => n7133, B => n6541, C => n7134, D => n6543, Z => 
                           n7132);
   U6737 : EO port map( A => n7135, B => n7136, Z => n7134);
   U6738 : EO port map( A => n6932, B => n7137, Z => n7136);
   U6739 : EN port map( A => n4921, B => n6969, Z => n7135);
   U6740 : EO port map( A => n7138, B => n7139, Z => n7133);
   U6741 : EO port map( A => n6939, B => n7140, Z => n7139);
   U6742 : EN port map( A => n5624, B => n6978, Z => n7138);
   U6743 : AO2 port map( A => n6440, B => n7141, C => n6551, D => n7142, Z => 
                           n7130);
   U6744 : EO port map( A => n7143, B => n7144, Z => n7142);
   U6745 : EO port map( A => n6946, B => n7145, Z => n7144);
   U6746 : EN port map( A => n4625, B => n6987, Z => n7143);
   U6747 : EO port map( A => v_KEY_COLUMN_28_port, B => v_DATA_COLUMN_28_port, 
                           Z => n7141);
   U6748 : EO port map( A => n7146, B => n7147, Z => n7129);
   U6749 : EO port map( A => n6953, B => n7148, Z => n7147);
   U6750 : EN port map( A => n4763, B => n6995, Z => n7146);
   U6751 : MUX21H port map( A => t_STATE_RAM0_0_28_port, B => v_RAM_IN0_28_port
                           , S => n6480, Z => n4064);
   U6752 : MUX21H port map( A => t_STATE_RAM0_1_28_port, B => v_RAM_IN0_28_port
                           , S => n6481, Z => n4063);
   U6753 : MUX21H port map( A => t_STATE_RAM0_2_28_port, B => v_RAM_IN0_28_port
                           , S => n6482, Z => n4062);
   U6754 : MUX21H port map( A => t_STATE_RAM0_3_28_port, B => v_RAM_IN0_28_port
                           , S => n4498, Z => n4061);
   U6755 : AO3 port map( A => n6483, B => n4447, C => n7149, D => n7150, Z => 
                           n4060);
   U6756 : AO2 port map( A => t_STATE_RAM0_3_28_port, B => n6486, C => 
                           v_RAM_OUT0_28_port, D => n4513, Z => n7150);
   U6757 : AO2 port map( A => t_STATE_RAM0_1_28_port, B => n4564, C => 
                           t_STATE_RAM0_2_28_port, D => n4563, Z => n7149);
   U6758 : AO3 port map( A => n7151, B => n6444, C => n7152, D => n7153, Z => 
                           n4059);
   U6759 : AO6 port map( A => v_RAM_IN0_12_port, B => n6538, C => n7154, Z => 
                           n7153);
   U6760 : AO4 port map( A => n7155, B => n6541, C => n7156, D => n6543, Z => 
                           n7154);
   U6761 : EO port map( A => n7157, B => n7158, Z => n7156);
   U6762 : EO port map( A => n6931, B => n7137, Z => n7158);
   U6763 : EO port map( A => n7159, B => n7160, Z => n7137);
   U6764 : EN port map( A => n6634, B => n6967, Z => n7160);
   U6765 : EN port map( A => n7161, B => n7162, Z => n6967);
   U6766 : EO port map( A => n6477, B => n7163, Z => n7161);
   U6767 : IV port map( A => n6820, Z => n6634);
   U6768 : EO port map( A => n4861, B => n4940, Z => n6820);
   U6769 : EN port map( A => n4958, B => n6970, Z => n7157);
   U6770 : IV port map( A => n6933, Z => n4958);
   U6771 : EO port map( A => n7164, B => n7165, Z => n7155);
   U6772 : EO port map( A => n6938, B => n7140, Z => n7165);
   U6773 : EO port map( A => n7166, B => n7167, Z => n7140);
   U6774 : EN port map( A => n6642, B => n6975, Z => n7167);
   U6775 : EN port map( A => n7168, B => n7169, Z => n6975);
   U6776 : EO port map( A => n6812, B => n7170, Z => n7168);
   U6777 : IV port map( A => n6813, Z => n6642);
   U6778 : EO port map( A => n5215, B => n6030, Z => n6813);
   U6779 : EO port map( A => n6490, B => n6979, Z => n7164);
   U6780 : AO2 port map( A => n6440, B => n7171, C => n6551, D => n7172, Z => 
                           n7152);
   U6781 : EO port map( A => n7173, B => n7174, Z => n7172);
   U6782 : EO port map( A => n6945, B => n7145, Z => n7174);
   U6783 : EN port map( A => n7175, B => n7176, Z => n7145);
   U6784 : EN port map( A => n6652, B => n6986, Z => n7176);
   U6785 : EN port map( A => n7177, B => n7178, Z => n6986);
   U6786 : EO port map( A => n6449, B => n7179, Z => n7177);
   U6787 : IV port map( A => n6796, Z => n6652);
   U6788 : EO port map( A => n4595, B => n4691, Z => n6796);
   U6789 : EN port map( A => n4718, B => n6988, Z => n7173);
   U6790 : IV port map( A => n6947, Z => n4718);
   U6791 : EO port map( A => v_KEY_COLUMN_12_port, B => v_DATA_COLUMN_12_port, 
                           Z => n7171);
   U6792 : EO port map( A => n7180, B => n7181, Z => n7151);
   U6793 : EO port map( A => n6952, B => n7148, Z => n7181);
   U6794 : EO port map( A => n7182, B => n7183, Z => n7148);
   U6795 : EN port map( A => n6660, B => n6993, Z => n7183);
   U6796 : EN port map( A => n7184, B => n7185, Z => n6993);
   U6797 : EO port map( A => n6461, B => n7186, Z => n7184);
   U6798 : IV port map( A => n6803, Z => n6660);
   U6799 : EO port map( A => n4743, B => n4784, Z => n6803);
   U6800 : EN port map( A => n4842, B => n6996, Z => n7180);
   U6801 : IV port map( A => n6954, Z => n4842);
   U6802 : MUX21H port map( A => t_STATE_RAM0_0_12_port, B => v_RAM_IN0_12_port
                           , S => n6480, Z => n4058);
   U6803 : MUX21H port map( A => t_STATE_RAM0_1_12_port, B => v_RAM_IN0_12_port
                           , S => n6481, Z => n4057);
   U6804 : MUX21H port map( A => t_STATE_RAM0_2_12_port, B => v_RAM_IN0_12_port
                           , S => n6482, Z => n4056);
   U6805 : MUX21H port map( A => t_STATE_RAM0_3_12_port, B => v_RAM_IN0_12_port
                           , S => n4498, Z => n4055);
   U6806 : AO3 port map( A => n6483, B => n4448, C => n7187, D => n7188, Z => 
                           n4054);
   U6807 : AO2 port map( A => t_STATE_RAM0_3_12_port, B => n6486, C => 
                           v_RAM_OUT0_12_port, D => n4513, Z => n7188);
   U6808 : AO2 port map( A => t_STATE_RAM0_1_12_port, B => n4564, C => 
                           t_STATE_RAM0_2_12_port, D => n4563, Z => n7187);
   U6809 : AO3 port map( A => n7189, B => n6444, C => n7190, D => n7191, Z => 
                           n4053);
   U6810 : AO6 port map( A => v_RAM_IN0_20_port, B => n6538, C => n7192, Z => 
                           n7191);
   U6811 : AO4 port map( A => n7193, B => n6541, C => n7194, D => n6543, Z => 
                           n7192);
   U6812 : EO port map( A => n7195, B => n7196, Z => n7194);
   U6813 : EO port map( A => n6932, B => n7197, Z => n7196);
   U6814 : EN port map( A => n7198, B => n4960, Z => n6932);
   U6815 : EN port map( A => n4861, B => n6970, Z => n7195);
   U6816 : EN port map( A => n7199, B => n4942, Z => n6970);
   U6817 : IV port map( A => n6965, Z => n4861);
   U6818 : EO port map( A => v_KEY_COLUMN_4_port, B => n7854, Z => n6965);
   U6819 : EO port map( A => n7200, B => n7201, Z => n7193);
   U6820 : EO port map( A => n6939, B => n7202, Z => n7201);
   U6821 : EO port map( A => n6229, B => n6664, Z => n6939);
   U6822 : EN port map( A => n5215, B => n6979, Z => n7200);
   U6823 : EO port map( A => n5821, B => n6076, Z => n6979);
   U6824 : IV port map( A => n6973, Z => n5215);
   U6825 : EO port map( A => v_KEY_COLUMN_4_port, B => n7920, Z => n6973);
   U6826 : AO2 port map( A => n6440, B => n7203, C => n6551, D => n7204, Z => 
                           n7190);
   U6827 : EO port map( A => n7205, B => n7206, Z => n7204);
   U6828 : EO port map( A => n6946, B => n7207, Z => n7206);
   U6829 : EN port map( A => n7208, B => n4721, Z => n6946);
   U6830 : EN port map( A => n4595, B => n6988, Z => n7205);
   U6831 : EN port map( A => n7209, B => n4694, Z => n6988);
   U6832 : IV port map( A => n6984, Z => n4595);
   U6833 : EO port map( A => v_KEY_COLUMN_4_port, B => n7852, Z => n6984);
   U6834 : EO port map( A => v_KEY_COLUMN_20_port, B => v_DATA_COLUMN_20_port, 
                           Z => n7203);
   U6835 : EO port map( A => n7210, B => n7211, Z => n7189);
   U6836 : EO port map( A => n6953, B => n7212, Z => n7211);
   U6837 : EN port map( A => n6457, B => n4844, Z => n6953);
   U6838 : EN port map( A => n4743, B => n6996, Z => n7210);
   U6839 : EN port map( A => n7213, B => n4786, Z => n6996);
   U6840 : IV port map( A => n6991, Z => n4743);
   U6841 : EO port map( A => v_KEY_COLUMN_4_port, B => n7917, Z => n6991);
   U6842 : MUX21H port map( A => t_STATE_RAM0_0_20_port, B => v_RAM_IN0_20_port
                           , S => n6480, Z => n4052);
   U6843 : MUX21H port map( A => t_STATE_RAM0_1_20_port, B => v_RAM_IN0_20_port
                           , S => n6481, Z => n4051);
   U6844 : MUX21H port map( A => t_STATE_RAM0_2_20_port, B => v_RAM_IN0_20_port
                           , S => n6482, Z => n4050);
   U6845 : MUX21H port map( A => t_STATE_RAM0_3_20_port, B => v_RAM_IN0_20_port
                           , S => n4498, Z => n4049);
   U6846 : AO3 port map( A => n6483, B => n4449, C => n7214, D => n7215, Z => 
                           n4048);
   U6847 : AO2 port map( A => t_STATE_RAM0_3_20_port, B => n6486, C => 
                           v_RAM_OUT0_20_port, D => n4513, Z => n7215);
   U6848 : AO2 port map( A => t_STATE_RAM0_1_20_port, B => n4564, C => 
                           t_STATE_RAM0_2_20_port, D => n4563, Z => n7214);
   U6849 : AO3 port map( A => n7216, B => n6444, C => n7217, D => n7218, Z => 
                           n4047);
   U6850 : AO6 port map( A => v_RAM_IN0_4_port, B => n6538, C => n7219, Z => 
                           n7218);
   U6851 : AO4 port map( A => n7220, B => n6541, C => n7221, D => n6543, Z => 
                           n7219);
   U6852 : EO port map( A => n7222, B => n7223, Z => n7221);
   U6853 : EO port map( A => n6931, B => n7197, Z => n7223);
   U6854 : EO port map( A => n7159, B => n7224, Z => n7197);
   U6855 : EN port map( A => n6633, B => n6968, Z => n7224);
   U6856 : EO port map( A => n7225, B => n7226, Z => n6968);
   U6857 : EO port map( A => n6782, B => n7227, Z => n7225);
   U6858 : EN port map( A => n4921, B => n6933, Z => n6633);
   U6859 : EO port map( A => v_KEY_COLUMN_28_port, B => n7856, Z => n6933);
   U6860 : EN port map( A => v_KEY_COLUMN_12_port, B => n7822, Z => n4921);
   U6861 : EN port map( A => n7228, B => n7229, Z => n7159);
   U6862 : EO port map( A => n7230, B => n7231, Z => n7229);
   U6863 : EO port map( A => n7232, B => n7233, Z => n7228);
   U6864 : EO port map( A => n6478, B => n7234, Z => n7233);
   U6865 : EN port map( A => n6635, B => n4923, Z => n6931);
   U6866 : EN port map( A => n4940, B => n6969, Z => n7222);
   U6867 : EN port map( A => n7235, B => n4863, Z => n6969);
   U6868 : EN port map( A => v_KEY_COLUMN_20_port, B => n7919, Z => n4940);
   U6869 : EO port map( A => n7236, B => n7237, Z => n7220);
   U6870 : EO port map( A => n6938, B => n7202, Z => n7237);
   U6871 : EO port map( A => n7166, B => n7238, Z => n7202);
   U6872 : EN port map( A => n6641, B => n6976, Z => n7238);
   U6873 : EO port map( A => n7239, B => n7240, Z => n6976);
   U6874 : EO port map( A => n6777, B => n7241, Z => n7239);
   U6875 : EN port map( A => n5624, B => n6490, Z => n6641);
   U6876 : EO port map( A => v_KEY_COLUMN_28_port, B => n7918, Z => n6490);
   U6877 : EN port map( A => v_KEY_COLUMN_12_port, B => n7812, Z => n5624);
   U6878 : EN port map( A => n7242, B => n7243, Z => n7166);
   U6879 : EO port map( A => n7244, B => n7245, Z => n7243);
   U6880 : EO port map( A => n7246, B => n7247, Z => n7242);
   U6881 : EO port map( A => n6468, B => n7248, Z => n7247);
   U6882 : EN port map( A => n6643, B => n5671, Z => n6938);
   U6883 : EN port map( A => n6030, B => n6978, Z => n7236);
   U6884 : EN port map( A => n6472, B => n5257, Z => n6978);
   U6885 : EN port map( A => v_KEY_COLUMN_20_port, B => n7807, Z => n6030);
   U6886 : AO2 port map( A => n6440, B => n7249, C => n6551, D => n7250, Z => 
                           n7217);
   U6887 : EO port map( A => n7251, B => n7252, Z => n7250);
   U6888 : EO port map( A => n6945, B => n7207, Z => n7252);
   U6889 : EN port map( A => n7175, B => n7253, Z => n7207);
   U6890 : EO port map( A => n6651, B => n6985, Z => n7253);
   U6891 : EN port map( A => n7254, B => n7255, Z => n6985);
   U6892 : EO port map( A => n6765, B => n7256, Z => n7254);
   U6893 : EN port map( A => n4625, B => n6947, Z => n6651);
   U6894 : EO port map( A => v_KEY_COLUMN_28_port, B => n7916, Z => n6947);
   U6895 : EN port map( A => v_KEY_COLUMN_12_port, B => n7846, Z => n4625);
   U6896 : EN port map( A => n7257, B => n7258, Z => n7175);
   U6897 : EN port map( A => n7259, B => n7260, Z => n7258);
   U6898 : EO port map( A => n7261, B => n7262, Z => n7257);
   U6899 : EO port map( A => n6451, B => n7263, Z => n7262);
   U6900 : EN port map( A => n6653, B => n4628, Z => n6945);
   U6901 : EN port map( A => n4691, B => n6987, Z => n7251);
   U6902 : EN port map( A => n7264, B => n4598, Z => n6987);
   U6903 : EN port map( A => v_KEY_COLUMN_20_port, B => n7915, Z => n4691);
   U6904 : EO port map( A => v_KEY_COLUMN_4_port, B => v_DATA_COLUMN_4_port, Z 
                           => n7249);
   U6905 : EO port map( A => n7265, B => n7266, Z => n7216);
   U6906 : EO port map( A => n6952, B => n7212, Z => n7266);
   U6907 : EO port map( A => n7182, B => n7267, Z => n7212);
   U6908 : EN port map( A => n6659, B => n6994, Z => n7267);
   U6909 : EO port map( A => n7268, B => n7269, Z => n6994);
   U6910 : EO port map( A => n6770, B => n7270, Z => n7268);
   U6911 : EN port map( A => n4763, B => n6954, Z => n6659);
   U6912 : EO port map( A => v_KEY_COLUMN_28_port, B => n7857, Z => n6954);
   U6913 : EN port map( A => v_KEY_COLUMN_12_port, B => n7841, Z => n4763);
   U6914 : EN port map( A => n7271, B => n7272, Z => n7182);
   U6915 : EO port map( A => n7273, B => n7274, Z => n7272);
   U6916 : EO port map( A => n7275, B => n7276, Z => n7271);
   U6917 : EO port map( A => n6458, B => n7277, Z => n7276);
   U6918 : EN port map( A => n6661, B => n4765, Z => n6952);
   U6919 : EN port map( A => n4784, B => n6995, Z => n7265);
   U6920 : EN port map( A => n7278, B => n4745, Z => n6995);
   U6921 : EN port map( A => v_KEY_COLUMN_20_port, B => n7834, Z => n4784);
   U6922 : MUX21H port map( A => t_STATE_RAM0_0_4_port, B => v_RAM_IN0_4_port, 
                           S => n6480, Z => n4046);
   U6923 : MUX21H port map( A => t_STATE_RAM0_1_4_port, B => v_RAM_IN0_4_port, 
                           S => n6481, Z => n4045);
   U6924 : MUX21H port map( A => t_STATE_RAM0_2_4_port, B => v_RAM_IN0_4_port, 
                           S => n6482, Z => n4044);
   U6925 : MUX21H port map( A => t_STATE_RAM0_3_4_port, B => v_RAM_IN0_4_port, 
                           S => n4498, Z => n4043);
   U6926 : AO3 port map( A => n6483, B => n4450, C => n7279, D => n7280, Z => 
                           n4042);
   U6927 : AO2 port map( A => t_STATE_RAM0_3_4_port, B => n6486, C => 
                           v_RAM_OUT0_4_port, D => n4513, Z => n7280);
   U6928 : AO2 port map( A => t_STATE_RAM0_1_4_port, B => n4564, C => 
                           t_STATE_RAM0_2_4_port, D => n4563, Z => n7279);
   U6929 : AO3 port map( A => n7281, B => n6444, C => n7282, D => n7283, Z => 
                           n4041);
   U6930 : AO6 port map( A => v_RAM_IN0_1_port, B => n6538, C => n7284, Z => 
                           n7283);
   U6931 : AO4 port map( A => n7285, B => n6541, C => n7286, D => n6543, Z => 
                           n7284);
   U6932 : EO port map( A => n7287, B => n7288, Z => n7286);
   U6933 : EN port map( A => n7107, B => n7289, Z => n7288);
   U6934 : EN port map( A => n4984, B => n7290, Z => n7287);
   U6935 : EO port map( A => n7291, B => n7292, Z => n7285);
   U6936 : EN port map( A => n7113, B => n7293, Z => n7292);
   U6937 : EN port map( A => n7294, B => n7029, Z => n7291);
   U6938 : AO2 port map( A => n6440, B => n7295, C => n6551, D => n7296, Z => 
                           n7282);
   U6939 : EO port map( A => n7297, B => n7298, Z => n7296);
   U6940 : EO port map( A => n7119, B => n7299, Z => n7298);
   U6941 : EN port map( A => n4727, B => n7300, Z => n7297);
   U6942 : EO port map( A => v_KEY_COLUMN_1_port, B => v_DATA_COLUMN_1_port, Z 
                           => n7295);
   U6943 : EO port map( A => n7301, B => n7302, Z => n7281);
   U6944 : EN port map( A => n7125, B => n7303, Z => n7302);
   U6945 : EN port map( A => n4848, B => n7304, Z => n7301);
   U6946 : MUX21H port map( A => t_STATE_RAM0_0_1_port, B => v_RAM_IN0_1_port, 
                           S => n6480, Z => n4040);
   U6947 : MUX21H port map( A => t_STATE_RAM0_1_1_port, B => v_RAM_IN0_1_port, 
                           S => n6481, Z => n4039);
   U6948 : MUX21H port map( A => t_STATE_RAM0_2_1_port, B => v_RAM_IN0_1_port, 
                           S => n6482, Z => n4038);
   U6949 : MUX21H port map( A => t_STATE_RAM0_3_1_port, B => v_RAM_IN0_1_port, 
                           S => n4498, Z => n4037);
   U6950 : AO3 port map( A => n6483, B => n4451, C => n7305, D => n7306, Z => 
                           n4036);
   U6951 : AO2 port map( A => t_STATE_RAM0_3_1_port, B => n6486, C => 
                           v_RAM_OUT0_1_port, D => n4513, Z => n7306);
   U6952 : AO2 port map( A => t_STATE_RAM0_1_1_port, B => n4564, C => 
                           t_STATE_RAM0_2_1_port, D => n4563, Z => n7305);
   U6953 : AO7 port map( A => n7307, B => n5009, C => n7308, Z => n4035);
   U6954 : AO2 port map( A => n6231, B => n4732, C => n7942, D => n6232, Z => 
                           n7308);
   U6955 : MUX21L port map( A => n7309, B => n7310, S => n4396, Z => n4732);
   U6956 : AO6 port map( A => v_RAM_OUT0_29_port, B => n7311, C => n4992, Z => 
                           n7310);
   U6957 : AO3 port map( A => n6278, B => n7312, C => n7313, D => n7314, Z => 
                           n4992);
   U6958 : ND4 port map( A => n7315, B => n7316, C => n7317, D => n7318, Z => 
                           n7314);
   U6959 : NR2 port map( A => v_RAM_OUT0_29_port, B => n7319, Z => n7318);
   U6960 : AO6 port map( A => n6293, B => n6505, C => n6337, Z => n7319);
   U6961 : IV port map( A => n6381, Z => n6505);
   U6962 : NR2 port map( A => v_RAM_OUT0_24_port, B => n6287, Z => n6381);
   U6963 : IV port map( A => n4996, Z => n6293);
   U6964 : AO2 port map( A => n6700, B => n6840, C => n6368, D => n6858, Z => 
                           n7317);
   U6965 : ND2 port map( A => n6506, B => n6341, Z => n6858);
   U6966 : IV port map( A => n6289, Z => n6341);
   U6967 : NR2 port map( A => n4355, B => n6287, Z => n6289);
   U6968 : ND2 port map( A => n4978, B => n6506, Z => n6840);
   U6969 : IV port map( A => n6837, Z => n4978);
   U6970 : AO2 port map( A => n6701, B => n6369, C => n6690, D => n6287, Z => 
                           n7316);
   U6971 : NR2 port map( A => n4355, B => n4413, Z => n6701);
   U6972 : AO2 port map( A => n6696, B => n6350, C => n6377, D => n4368, Z => 
                           n7315);
   U6973 : ND3 port map( A => n6519, B => n7320, C => n7321, Z => n7313);
   U6974 : AO1 port map( A => n4996, B => n6265, C => n6277, D => n7322, Z => 
                           n7321);
   U6975 : NR2 port map( A => n6346, B => n6326, Z => n7322);
   U6976 : NR2 port map( A => n6688, B => n4355, Z => n6346);
   U6977 : IV port map( A => n6712, Z => n6688);
   U6978 : NR2 port map( A => v_RAM_OUT0_27_port, B => v_RAM_OUT0_24_port, Z =>
                           n6277);
   U6979 : AO4 port map( A => n6253, B => n6301, C => n4975, D => n7323, Z => 
                           n7320);
   U6980 : NR2 port map( A => v_RAM_OUT0_28_port, B => n6427, Z => n7323);
   U6981 : IV port map( A => n6301, Z => n6427);
   U6982 : NR2 port map( A => v_RAM_OUT0_24_port, B => n6712, Z => n6301);
   U6983 : NR2 port map( A => n4404, B => v_RAM_OUT0_25_port, Z => n6519);
   U6984 : ND2 port map( A => n4994, B => n5004, Z => n7312);
   U6985 : IV port map( A => n4993, Z => n5004);
   U6986 : NR2 port map( A => n4364, B => n4404, Z => n4994);
   U6987 : IV port map( A => n7324, Z => n6278);
   U6988 : AO4 port map( A => n4996, B => n6300, C => n6311, D => n4997, Z => 
                           n7311);
   U6989 : IV port map( A => n6432, Z => n4997);
   U6990 : NR2 port map( A => n6239, B => n6299, Z => n6432);
   U6991 : NR2 port map( A => n4976, B => v_RAM_OUT0_24_port, Z => n6299);
   U6992 : IV port map( A => n6700, Z => n6311);
   U6993 : IV port map( A => n6368, Z => n6300);
   U6994 : NR2 port map( A => n6326, B => n4364, Z => n6368);
   U6995 : AO3 port map( A => n6398, B => n6240, C => n7325, D => n7326, Z => 
                           n7309);
   U6996 : AO2 port map( A => n6250, B => n5000, C => v_RAM_OUT0_29_port, D => 
                           n5007, Z => n7326);
   U6997 : ND4 port map( A => n7327, B => n7328, C => n7329, D => n7330, Z => 
                           n5007);
   U6998 : AO2 port map( A => v_RAM_OUT0_25_port, B => n7331, C => n6510, D => 
                           n6690, Z => n7330);
   U6999 : NR2 port map( A => n4979, B => v_RAM_OUT0_25_port, Z => n6690);
   U7000 : AO4 port map( A => n4410, B => n6291, C => n7332, D => n4359, Z => 
                           n7331);
   U7001 : NR2 port map( A => n6308, B => n6367, Z => n7332);
   U7002 : ND2 port map( A => n4355, B => n6340, Z => n6291);
   U7003 : AO2 port map( A => n6365, B => n6284, C => n6359, D => n7049, Z => 
                           n7329);
   U7004 : IV port map( A => n6428, Z => n7049);
   U7005 : NR2 port map( A => n6290, B => n6846, Z => n6428);
   U7006 : NR2 port map( A => n6337, B => n4364, Z => n6359);
   U7007 : ND2 port map( A => n6506, B => n6314, Z => n6284);
   U7008 : IV port map( A => n6367, Z => n6314);
   U7009 : NR2 port map( A => n4355, B => n6403, Z => n6367);
   U7010 : IV port map( A => n6288, Z => n6403);
   U7011 : NR2 port map( A => n6337, B => v_RAM_OUT0_25_port, Z => n6365);
   U7012 : AO2 port map( A => n6700, B => n6350, C => n6837, D => n6369, Z => 
                           n7328);
   U7013 : NR2 port map( A => n4979, B => n4364, Z => n6369);
   U7014 : IV port map( A => n6333, Z => n4979);
   U7015 : NR2 port map( A => n4355, B => n6712, Z => n6837);
   U7016 : ND2 port map( A => v_RAM_OUT0_24_port, B => n4976, Z => n6350);
   U7017 : IV port map( A => n6330, Z => n4976);
   U7018 : NR2 port map( A => n4364, B => n6329, Z => n6700);
   U7019 : AO2 port map( A => n6377, B => n6330, C => n6696, D => n6370, Z => 
                           n7327);
   U7020 : ND2 port map( A => n6410, B => n4980, Z => n6370);
   U7021 : IV port map( A => n6846, Z => n4980);
   U7022 : NR2 port map( A => v_RAM_OUT0_30_port, B => v_RAM_OUT0_24_port, Z =>
                           n6846);
   U7023 : IV port map( A => n6239, Z => n6410);
   U7024 : NR2 port map( A => n6340, B => n4355, Z => n6239);
   U7025 : NR2 port map( A => n6329, B => v_RAM_OUT0_25_port, Z => n6696);
   U7026 : NR2 port map( A => n6326, B => v_RAM_OUT0_25_port, Z => n6377);
   U7027 : AO7 port map( A => n6521, B => n6337, C => n7333, Z => n5000);
   U7028 : AO2 port map( A => n7324, B => n7334, C => n6510, D => n4975, Z => 
                           n7333);
   U7029 : NR2 port map( A => n4996, B => n6712, Z => n6510);
   U7030 : AO7 port map( A => n4359, B => n6339, C => n6326, Z => n7334);
   U7031 : IV port map( A => n6308, Z => n6339);
   U7032 : NR2 port map( A => n6352, B => v_RAM_OUT0_24_port, Z => n6308);
   U7033 : IV port map( A => n6287, Z => n6352);
   U7034 : NR2 port map( A => n6253, B => n4967, Z => n7324);
   U7035 : NR2 port map( A => n4355, B => v_RAM_OUT0_27_port, Z => n6253);
   U7036 : IV port map( A => n6265, Z => n6337);
   U7037 : NR2 port map( A => n6290, B => n6426, Z => n6521);
   U7038 : NR2 port map( A => n6340, B => v_RAM_OUT0_24_port, Z => n6426);
   U7039 : IV port map( A => n6347, Z => n6340);
   U7040 : NR2 port map( A => n4368, B => n4355, Z => n6290);
   U7041 : NR2 port map( A => v_RAM_OUT0_29_port, B => v_RAM_OUT0_25_port, Z =>
                           n6250);
   U7042 : AO2 port map( A => n7335, B => n6252, C => n5005, D => n6254, Z => 
                           n7325);
   U7043 : NR2 port map( A => n4982, B => n6326, Z => n6254);
   U7044 : IV port map( A => n6281, Z => n6326);
   U7045 : NR2 port map( A => n4359, B => v_RAM_OUT0_28_port, Z => n6281);
   U7046 : NR2 port map( A => n6288, B => n4996, Z => n5005);
   U7047 : NR2 port map( A => n4355, B => n6347, Z => n4996);
   U7048 : NR2 port map( A => n4413, B => v_RAM_OUT0_27_port, Z => n6288);
   U7049 : NR2 port map( A => n5003, B => n4993, Z => n7335);
   U7050 : NR2 port map( A => n6333, B => n6265, Z => n4993);
   U7051 : NR2 port map( A => v_RAM_OUT0_28_port, B => v_RAM_OUT0_26_port, Z =>
                           n6265);
   U7052 : NR2 port map( A => n4359, B => n4410, Z => n6333);
   U7053 : IV port map( A => n6709, Z => n5003);
   U7054 : ND2 port map( A => n6506, B => n6275, Z => n6709);
   U7055 : ND2 port map( A => n6287, B => v_RAM_OUT0_24_port, Z => n6275);
   U7056 : NR2 port map( A => n4368, B => v_RAM_OUT0_30_port, Z => n6287);
   U7057 : ND2 port map( A => v_RAM_OUT0_30_port, B => n4355, Z => n6506);
   U7058 : IV port map( A => n6292, Z => n6240);
   U7059 : NR2 port map( A => n4982, B => n6329, Z => n6292);
   U7060 : IV port map( A => n4975, Z => n6329);
   U7061 : NR2 port map( A => n4410, B => v_RAM_OUT0_26_port, Z => n4975);
   U7062 : IV port map( A => n6252, Z => n4982);
   U7063 : NR2 port map( A => n4364, B => v_RAM_OUT0_29_port, Z => n6252);
   U7064 : NR2 port map( A => n4967, B => n6276, Z => n6398);
   U7065 : NR2 port map( A => n4355, B => v_RAM_OUT0_30_port, Z => n6276);
   U7066 : NR2 port map( A => v_RAM_OUT0_24_port, B => n6330, Z => n4967);
   U7067 : NR2 port map( A => n6347, B => n6712, Z => n6330);
   U7068 : NR2 port map( A => n4368, B => n4413, Z => n6712);
   U7069 : NR2 port map( A => v_RAM_OUT0_30_port, B => v_RAM_OUT0_27_port, Z =>
                           n6347);
   U7070 : NR2 port map( A => n5384, B => n6232, Z => n6231);
   U7071 : NR2 port map( A => n5384, B => n4611, Z => n6232);
   U7072 : AN3 port map( A => n4560, B => n4399, C => n6228, Z => n4611);
   U7073 : NR2 port map( A => v_CALCULATION_CNTR_3_port, B => 
                           v_CALCULATION_CNTR_2_port, Z => n4560);
   U7074 : AO3 port map( A => n7336, B => n6444, C => n7337, D => n7338, Z => 
                           n4034);
   U7075 : AO6 port map( A => v_RAM_IN0_25_port, B => n6538, C => n7339, Z => 
                           n7338);
   U7076 : AO4 port map( A => n7340, B => n6541, C => n7341, D => n6543, Z => 
                           n7339);
   U7077 : EO port map( A => n7342, B => n7343, Z => n7341);
   U7078 : EO port map( A => n7289, B => n7344, Z => n7343);
   U7079 : EN port map( A => n7345, B => n7346, Z => n7289);
   U7080 : EO port map( A => n6479, B => n7347, Z => n7346);
   U7081 : EN port map( A => n4888, B => n7109, Z => n7342);
   U7082 : EO port map( A => n7348, B => n7349, Z => n7340);
   U7083 : EO port map( A => n7293, B => n7350, Z => n7349);
   U7084 : EN port map( A => n7351, B => n7352, Z => n7293);
   U7085 : EO port map( A => n7082, B => n7353, Z => n7352);
   U7086 : EN port map( A => n5345, B => n7114, Z => n7348);
   U7087 : AO2 port map( A => n6440, B => n7354, C => n6551, D => n7355, Z => 
                           n7337);
   U7088 : EO port map( A => n7356, B => n7357, Z => n7355);
   U7089 : EN port map( A => n7299, B => n7358, Z => n7357);
   U7090 : EN port map( A => n7359, B => n7360, Z => n7299);
   U7091 : EO port map( A => n6453, B => n7361, Z => n7360);
   U7092 : EN port map( A => n4604, B => n7121, Z => n7356);
   U7093 : EO port map( A => v_KEY_COLUMN_25_port, B => v_DATA_COLUMN_25_port, 
                           Z => n7354);
   U7094 : EO port map( A => n7362, B => n7363, Z => n7336);
   U7095 : EO port map( A => n7303, B => n7364, Z => n7363);
   U7096 : EN port map( A => n7365, B => n7366, Z => n7303);
   U7097 : EO port map( A => n6456, B => n7367, Z => n7366);
   U7098 : EN port map( A => n4749, B => n7126, Z => n7362);
   U7099 : MUX21H port map( A => t_STATE_RAM0_0_25_port, B => v_RAM_IN0_25_port
                           , S => n6480, Z => n4033);
   U7100 : MUX21H port map( A => t_STATE_RAM0_1_25_port, B => v_RAM_IN0_25_port
                           , S => n6481, Z => n4032);
   U7101 : MUX21H port map( A => t_STATE_RAM0_2_25_port, B => v_RAM_IN0_25_port
                           , S => n6482, Z => n4031);
   U7102 : MUX21H port map( A => t_STATE_RAM0_3_25_port, B => v_RAM_IN0_25_port
                           , S => n4498, Z => n4030);
   U7103 : AO3 port map( A => n6483, B => n4452, C => n7368, D => n7369, Z => 
                           n4029);
   U7104 : AO2 port map( A => t_STATE_RAM0_3_25_port, B => n6486, C => 
                           v_RAM_OUT0_25_port, D => n4513, Z => n7369);
   U7105 : AO2 port map( A => t_STATE_RAM0_1_25_port, B => n4564, C => 
                           t_STATE_RAM0_2_25_port, D => n4563, Z => n7368);
   U7106 : AO3 port map( A => n7370, B => n6444, C => n7371, D => n7372, Z => 
                           n4028);
   U7107 : AO6 port map( A => v_RAM_IN0_17_port, B => n6538, C => n7373, Z => 
                           n7372);
   U7108 : AO4 port map( A => n7374, B => n6541, C => n7375, D => n6543, Z => 
                           n7373);
   U7109 : EO port map( A => n7376, B => n7377, Z => n7375);
   U7110 : EO port map( A => n7108, B => n7344, Z => n7377);
   U7111 : EN port map( A => n7378, B => n7379, Z => n7108);
   U7112 : EO port map( A => n7073, B => n7347, Z => n7379);
   U7113 : EO port map( A => n6585, B => n7380, Z => n7347);
   U7114 : EO port map( A => n6477, B => n6546, Z => n7380);
   U7115 : EN port map( A => n6600, B => n7381, Z => n6546);
   U7116 : EN port map( A => n6930, B => n4935, Z => n6585);
   U7117 : IV port map( A => n6630, Z => n6930);
   U7118 : EN port map( A => n4927, B => n7290, Z => n7376);
   U7119 : EO port map( A => n7382, B => n7383, Z => n7374);
   U7120 : EO port map( A => n7112, B => n7350, Z => n7383);
   U7121 : EN port map( A => n7384, B => n7385, Z => n7112);
   U7122 : EO port map( A => n7081, B => n7353, Z => n7385);
   U7123 : EO port map( A => n6579, B => n7386, Z => n7353);
   U7124 : EN port map( A => n6812, B => n6547, Z => n7386);
   U7125 : EO port map( A => n6605, B => n5095, Z => n6547);
   U7126 : EN port map( A => n6937, B => n5907, Z => n6579);
   U7127 : EN port map( A => n5756, B => n7294, Z => n7382);
   U7128 : AO2 port map( A => n6440, B => n7387, C => n6551, D => n7388, Z => 
                           n7371);
   U7129 : EO port map( A => n7389, B => n7390, Z => n7388);
   U7130 : EN port map( A => n7120, B => n7358, Z => n7390);
   U7131 : EN port map( A => n7391, B => n7392, Z => n7120);
   U7132 : EO port map( A => n7088, B => n7361, Z => n7392);
   U7133 : EO port map( A => n6567, B => n7393, Z => n7361);
   U7134 : EN port map( A => n6449, B => n6555, Z => n7393);
   U7135 : EN port map( A => n6612, B => n4589, Z => n6555);
   U7136 : IV port map( A => n7394, Z => n4589);
   U7137 : EN port map( A => n7395, B => n4684, Z => n6567);
   U7138 : IV port map( A => n6648, Z => n7395);
   U7139 : EN port map( A => n4652, B => n7300, Z => n7389);
   U7140 : EO port map( A => v_KEY_COLUMN_17_port, B => v_DATA_COLUMN_17_port, 
                           Z => n7387);
   U7141 : EO port map( A => n7396, B => n7397, Z => n7370);
   U7142 : EO port map( A => n7124, B => n7364, Z => n7397);
   U7143 : EN port map( A => n7398, B => n7399, Z => n7124);
   U7144 : EO port map( A => n7094, B => n7367, Z => n7399);
   U7145 : EO port map( A => n6572, B => n7400, Z => n7367);
   U7146 : EN port map( A => n6461, B => n6556, Z => n7400);
   U7147 : EO port map( A => n6617, B => n7401, Z => n6556);
   U7148 : EN port map( A => n6951, B => n4779, Z => n6572);
   U7149 : IV port map( A => n6656, Z => n6951);
   U7150 : EN port map( A => n4770, B => n7304, Z => n7396);
   U7151 : MUX21H port map( A => t_STATE_RAM0_0_17_port, B => v_RAM_IN0_17_port
                           , S => n6480, Z => n4027);
   U7152 : MUX21H port map( A => t_STATE_RAM0_1_17_port, B => v_RAM_IN0_17_port
                           , S => n6481, Z => n4026);
   U7153 : MUX21H port map( A => t_STATE_RAM0_2_17_port, B => v_RAM_IN0_17_port
                           , S => n6482, Z => n4025);
   U7154 : MUX21H port map( A => t_STATE_RAM0_3_17_port, B => v_RAM_IN0_17_port
                           , S => n4498, Z => n4024);
   U7155 : AO3 port map( A => n6483, B => n4453, C => n7402, D => n7403, Z => 
                           n4023);
   U7156 : AO2 port map( A => t_STATE_RAM0_3_17_port, B => n6486, C => 
                           v_RAM_OUT0_17_port, D => n4513, Z => n7403);
   U7157 : AO2 port map( A => t_STATE_RAM0_1_17_port, B => n4564, C => 
                           t_STATE_RAM0_2_17_port, D => n4563, Z => n7402);
   U7158 : AO3 port map( A => n7404, B => n6444, C => n7405, D => n7406, Z => 
                           n4022);
   U7159 : AO6 port map( A => v_RAM_IN0_26_port, B => n6538, C => n7407, Z => 
                           n7406);
   U7160 : AO4 port map( A => n7408, B => n6541, C => n7409, D => n6543, Z => 
                           n7407);
   U7161 : EO port map( A => n7410, B => n7411, Z => n7409);
   U7162 : EN port map( A => n7412, B => n7378, Z => n7411);
   U7163 : EO port map( A => n4888, B => n4984, Z => n7378);
   U7164 : EN port map( A => n4944, B => n7072, Z => n7410);
   U7165 : EN port map( A => n7413, B => n7414, Z => n7072);
   U7166 : EN port map( A => n4865, B => n4925, Z => n7414);
   U7167 : EO port map( A => n7415, B => n7416, Z => n7408);
   U7168 : EN port map( A => n7417, B => n7384, Z => n7416);
   U7169 : EO port map( A => n5345, B => n7029, Z => n7384);
   U7170 : EN port map( A => n6125, B => n7078, Z => n7415);
   U7171 : EN port map( A => n7418, B => n7419, Z => n7078);
   U7172 : EN port map( A => n5305, B => n5713, Z => n7419);
   U7173 : AO2 port map( A => n6440, B => n7420, C => n6551, D => n7421, Z => 
                           n7405);
   U7174 : EO port map( A => n7422, B => n7423, Z => n7421);
   U7175 : EO port map( A => n7391, B => n7424, Z => n7423);
   U7176 : EO port map( A => n4604, B => n4727, Z => n7391);
   U7177 : EN port map( A => n4697, B => n7087, Z => n7422);
   U7178 : EN port map( A => n7425, B => n7426, Z => n7087);
   U7179 : EN port map( A => n4601, B => n4631, Z => n7426);
   U7180 : EO port map( A => v_KEY_COLUMN_26_port, B => v_DATA_COLUMN_26_port, 
                           Z => n7420);
   U7181 : EO port map( A => n7427, B => n7428, Z => n7404);
   U7182 : EN port map( A => n7429, B => n7398, Z => n7428);
   U7183 : EN port map( A => n4749, B => n7430, Z => n7398);
   U7184 : EN port map( A => n4788, B => n7093, Z => n7427);
   U7185 : EN port map( A => n7431, B => n7432, Z => n7093);
   U7186 : EN port map( A => n4747, B => n4767, Z => n7432);
   U7187 : MUX21H port map( A => t_STATE_RAM0_0_26_port, B => v_RAM_IN0_26_port
                           , S => n6480, Z => n4021);
   U7188 : MUX21H port map( A => t_STATE_RAM0_1_26_port, B => v_RAM_IN0_26_port
                           , S => n6481, Z => n4020);
   U7189 : MUX21H port map( A => t_STATE_RAM0_2_26_port, B => v_RAM_IN0_26_port
                           , S => n6482, Z => n4019);
   U7190 : MUX21H port map( A => t_STATE_RAM0_3_26_port, B => v_RAM_IN0_26_port
                           , S => n4498, Z => n4018);
   U7191 : AO3 port map( A => n6483, B => n4454, C => n7433, D => n7434, Z => 
                           n4017);
   U7192 : AO2 port map( A => t_STATE_RAM0_3_26_port, B => n6486, C => 
                           v_RAM_OUT0_26_port, D => n4513, Z => n7434);
   U7193 : AO2 port map( A => t_STATE_RAM0_1_26_port, B => n4564, C => 
                           t_STATE_RAM0_2_26_port, D => n4563, Z => n7433);
   U7194 : AO3 port map( A => n7435, B => n6444, C => n7436, D => n7437, Z => 
                           n4016);
   U7195 : AO6 port map( A => v_RAM_IN0_10_port, B => n6538, C => n7438, Z => 
                           n7437);
   U7196 : AO4 port map( A => n7439, B => n6541, C => n7440, D => n6543, Z => 
                           n7438);
   U7197 : EO port map( A => n7441, B => n7442, Z => n7440);
   U7198 : EN port map( A => n7412, B => n7345, Z => n7442);
   U7199 : EN port map( A => n4927, B => n7443, Z => n7345);
   U7200 : EN port map( A => n7107, B => n7344, Z => n7412);
   U7201 : EN port map( A => n4865, B => n7008, Z => n7441);
   U7202 : EN port map( A => n7413, B => n7444, Z => n7008);
   U7203 : EN port map( A => n4944, B => n4962, Z => n7444);
   U7204 : IV port map( A => n7075, Z => n4962);
   U7205 : EO port map( A => n7109, B => n7290, Z => n7413);
   U7206 : EN port map( A => n6782, B => n7445, Z => n7290);
   U7207 : EN port map( A => n4852, B => n4931, Z => n7445);
   U7208 : EN port map( A => n7446, B => n7447, Z => n7109);
   U7209 : EN port map( A => n4950, B => n4954, Z => n7447);
   U7210 : EN port map( A => n4912, B => n4918, Z => n7446);
   U7211 : EO port map( A => n7448, B => n7449, Z => n7439);
   U7212 : EN port map( A => n7417, B => n7351, Z => n7449);
   U7213 : EO port map( A => n5756, B => n6164, Z => n7351);
   U7214 : IV port map( A => n7450, Z => n5756);
   U7215 : EN port map( A => n7113, B => n7350, Z => n7417);
   U7216 : EN port map( A => n5305, B => n7013, Z => n7448);
   U7217 : EN port map( A => n7418, B => n7451, Z => n7013);
   U7218 : EN port map( A => n6125, B => n6826, Z => n7451);
   U7219 : IV port map( A => n7080, Z => n6826);
   U7220 : EO port map( A => n7294, B => n7114, Z => n7418);
   U7221 : EN port map( A => n7452, B => n7453, Z => n7114);
   U7222 : EN port map( A => n6229, B => n6315, Z => n7453);
   U7223 : IV port map( A => n6584, Z => n6315);
   U7224 : EN port map( A => n6643, B => n5507, Z => n7452);
   U7225 : EN port map( A => n6777, B => n7454, Z => n7294);
   U7226 : EN port map( A => n5008, B => n5821, Z => n7454);
   U7227 : AO2 port map( A => n6440, B => n7455, C => n6551, D => n7456, Z => 
                           n7436);
   U7228 : EO port map( A => n7457, B => n7458, Z => n7456);
   U7229 : EO port map( A => n7359, B => n7424, Z => n7458);
   U7230 : EN port map( A => n7119, B => n7358, Z => n7424);
   U7231 : IV port map( A => n7459, Z => n7358);
   U7232 : EN port map( A => n7460, B => n4700, Z => n7359);
   U7233 : EN port map( A => n4601, B => n7020, Z => n7457);
   U7234 : EN port map( A => n7425, B => n7461, Z => n7020);
   U7235 : EN port map( A => n4697, B => n4724, Z => n7461);
   U7236 : IV port map( A => n7090, Z => n4724);
   U7237 : EO port map( A => n7121, B => n7300, Z => n7425);
   U7238 : EN port map( A => n6765, B => n7462, Z => n7300);
   U7239 : EN port map( A => n4583, B => n4679, Z => n7462);
   U7240 : EN port map( A => n7463, B => n7464, Z => n7121);
   U7241 : EN port map( A => n4707, B => n4712, Z => n7464);
   U7242 : EN port map( A => n4613, B => n4621, Z => n7463);
   U7243 : EO port map( A => v_KEY_COLUMN_10_port, B => v_DATA_COLUMN_10_port, 
                           Z => n7455);
   U7244 : EO port map( A => n7465, B => n7466, Z => n7435);
   U7245 : EN port map( A => n7429, B => n7365, Z => n7466);
   U7246 : EN port map( A => n4770, B => n7467, Z => n7365);
   U7247 : EN port map( A => n7125, B => n7364, Z => n7429);
   U7248 : EN port map( A => n4747, B => n7025, Z => n7465);
   U7249 : EN port map( A => n7431, B => n7468, Z => n7025);
   U7250 : EN port map( A => n4788, B => n4846, Z => n7468);
   U7251 : IV port map( A => n7096, Z => n4846);
   U7252 : EO port map( A => n7126, B => n7304, Z => n7431);
   U7253 : EN port map( A => n6770, B => n7469, Z => n7304);
   U7254 : EN port map( A => n4734, B => n4775, Z => n7469);
   U7255 : EN port map( A => n7470, B => n7471, Z => n7126);
   U7256 : EN port map( A => n4834, B => n4838, Z => n7471);
   U7257 : EN port map( A => n4754, B => n4760, Z => n7470);
   U7258 : MUX21H port map( A => t_STATE_RAM0_0_10_port, B => v_RAM_IN0_10_port
                           , S => n6480, Z => n4015);
   U7259 : MUX21H port map( A => t_STATE_RAM0_1_10_port, B => v_RAM_IN0_10_port
                           , S => n6481, Z => n4014);
   U7260 : MUX21H port map( A => t_STATE_RAM0_2_10_port, B => v_RAM_IN0_10_port
                           , S => n6482, Z => n4013);
   U7261 : MUX21H port map( A => t_STATE_RAM0_3_10_port, B => v_RAM_IN0_10_port
                           , S => n4498, Z => n4012);
   U7262 : AO3 port map( A => n6483, B => n4455, C => n7472, D => n7473, Z => 
                           n4011);
   U7263 : AO2 port map( A => t_STATE_RAM0_3_10_port, B => n6486, C => 
                           v_RAM_OUT0_10_port, D => n4513, Z => n7473);
   U7264 : AO2 port map( A => t_STATE_RAM0_1_10_port, B => n4564, C => 
                           t_STATE_RAM0_2_10_port, D => n4563, Z => n7472);
   U7265 : AO3 port map( A => n7474, B => n6444, C => n7475, D => n7476, Z => 
                           n4010);
   U7266 : AO6 port map( A => v_RAM_IN0_27_port, B => n6538, C => n7477, Z => 
                           n7476);
   U7267 : AO4 port map( A => n7478, B => n6541, C => n7479, D => n6543, Z => 
                           n7477);
   U7268 : EO port map( A => n7480, B => n7481, Z => n7479);
   U7269 : EN port map( A => n7482, B => n7483, Z => n7481);
   U7270 : EO port map( A => n7162, B => n7484, Z => n7480);
   U7271 : EN port map( A => n4942, B => n7227, Z => n7484);
   U7272 : EO port map( A => n7485, B => n7486, Z => n7478);
   U7273 : EN port map( A => n7487, B => n7488, Z => n7486);
   U7274 : EO port map( A => n7169, B => n7489, Z => n7485);
   U7275 : EN port map( A => n6076, B => n7240, Z => n7489);
   U7276 : AO2 port map( A => n6440, B => n7490, C => n6551, D => n7491, Z => 
                           n7475);
   U7277 : EO port map( A => n7492, B => n7493, Z => n7491);
   U7278 : EO port map( A => n7494, B => n7495, Z => n7493);
   U7279 : EO port map( A => n7178, B => n7496, Z => n7492);
   U7280 : EN port map( A => n4694, B => n7256, Z => n7496);
   U7281 : EO port map( A => v_KEY_COLUMN_27_port, B => v_DATA_COLUMN_27_port, 
                           Z => n7490);
   U7282 : EO port map( A => n7497, B => n7498, Z => n7474);
   U7283 : EN port map( A => n7499, B => n7500, Z => n7498);
   U7284 : EO port map( A => n7185, B => n7501, Z => n7497);
   U7285 : EN port map( A => n4786, B => n7270, Z => n7501);
   U7286 : MUX21H port map( A => t_STATE_RAM0_0_27_port, B => v_RAM_IN0_27_port
                           , S => n6480, Z => n4009);
   U7287 : MUX21H port map( A => t_STATE_RAM0_1_27_port, B => v_RAM_IN0_27_port
                           , S => n6481, Z => n4008);
   U7288 : MUX21H port map( A => t_STATE_RAM0_2_27_port, B => v_RAM_IN0_27_port
                           , S => n6482, Z => n4007);
   U7289 : MUX21H port map( A => t_STATE_RAM0_3_27_port, B => v_RAM_IN0_27_port
                           , S => n4498, Z => n4006);
   U7290 : AO3 port map( A => n6483, B => n4456, C => n7502, D => n7503, Z => 
                           n4005);
   U7291 : AO2 port map( A => t_STATE_RAM0_3_27_port, B => n6486, C => 
                           v_RAM_OUT0_27_port, D => n4513, Z => n7503);
   U7292 : AO2 port map( A => t_STATE_RAM0_1_27_port, B => n4564, C => 
                           t_STATE_RAM0_2_27_port, D => n4563, Z => n7502);
   U7293 : AO3 port map( A => n7504, B => n6444, C => n7505, D => n7506, Z => 
                           n4004);
   U7294 : AO6 port map( A => v_RAM_IN0_19_port, B => n6538, C => n7507, Z => 
                           n7506);
   U7295 : AO4 port map( A => n7508, B => n6541, C => n7509, D => n6543, Z => 
                           n7507);
   U7296 : EO port map( A => n7510, B => n7511, Z => n7509);
   U7297 : EN port map( A => n7482, B => n7512, Z => n7511);
   U7298 : EN port map( A => n7513, B => n7514, Z => n7482);
   U7299 : EN port map( A => n4863, B => n4923, Z => n7514);
   U7300 : EO port map( A => n7162, B => n7515, Z => n7510);
   U7301 : EN port map( A => n4960, B => n7226, Z => n7515);
   U7302 : EN port map( A => n4950, B => n7075, Z => n7162);
   U7303 : EO port map( A => v_KEY_COLUMN_26_port, B => n7869, Z => n7075);
   U7304 : EO port map( A => n7516, B => n7517, Z => n7508);
   U7305 : EN port map( A => n7487, B => n7518, Z => n7517);
   U7306 : EN port map( A => n7519, B => n7520, Z => n7487);
   U7307 : EN port map( A => n5257, B => n5671, Z => n7520);
   U7308 : EO port map( A => n7169, B => n7521, Z => n7516);
   U7309 : EN port map( A => n6664, B => n7241, Z => n7521);
   U7310 : EN port map( A => n6229, B => n7080, Z => n7169);
   U7311 : EO port map( A => v_KEY_COLUMN_26_port, B => n7930, Z => n7080);
   U7312 : AO2 port map( A => n6440, B => n7522, C => n6551, D => n7523, Z => 
                           n7505);
   U7313 : EO port map( A => n7524, B => n7525, Z => n7523);
   U7314 : EO port map( A => n7494, B => n7526, Z => n7525);
   U7315 : EN port map( A => n7527, B => n7528, Z => n7494);
   U7316 : EN port map( A => n4598, B => n4628, Z => n7528);
   U7317 : EO port map( A => n7178, B => n7529, Z => n7524);
   U7318 : EN port map( A => n4721, B => n7255, Z => n7529);
   U7319 : EN port map( A => n4707, B => n7090, Z => n7178);
   U7320 : EO port map( A => v_KEY_COLUMN_26_port, B => n7928, Z => n7090);
   U7321 : EO port map( A => v_KEY_COLUMN_19_port, B => v_DATA_COLUMN_19_port, 
                           Z => n7522);
   U7322 : EO port map( A => n7530, B => n7531, Z => n7504);
   U7323 : EN port map( A => n7499, B => n7532, Z => n7531);
   U7324 : EN port map( A => n7533, B => n7534, Z => n7499);
   U7325 : EN port map( A => n4745, B => n4765, Z => n7534);
   U7326 : EO port map( A => n7185, B => n7535, Z => n7530);
   U7327 : EN port map( A => n4844, B => n7269, Z => n7535);
   U7328 : EN port map( A => n4834, B => n7096, Z => n7185);
   U7329 : EO port map( A => v_KEY_COLUMN_26_port, B => n7871, Z => n7096);
   U7330 : MUX21H port map( A => t_STATE_RAM0_0_19_port, B => v_RAM_IN0_19_port
                           , S => n6480, Z => n4003);
   U7331 : MUX21H port map( A => t_STATE_RAM0_1_19_port, B => v_RAM_IN0_19_port
                           , S => n6481, Z => n4002);
   U7332 : MUX21H port map( A => t_STATE_RAM0_2_19_port, B => v_RAM_IN0_19_port
                           , S => n6482, Z => n4001);
   U7333 : MUX21H port map( A => t_STATE_RAM0_3_19_port, B => v_RAM_IN0_19_port
                           , S => n4498, Z => n4000);
   U7334 : AO3 port map( A => n6483, B => n4457, C => n7536, D => n7537, Z => 
                           n3999);
   U7335 : AO2 port map( A => t_STATE_RAM0_3_19_port, B => n6486, C => 
                           v_RAM_OUT0_19_port, D => n4513, Z => n7537);
   U7336 : AO2 port map( A => t_STATE_RAM0_1_19_port, B => n4564, C => 
                           t_STATE_RAM0_2_19_port, D => n4563, Z => n7536);
   U7337 : AO3 port map( A => n7538, B => n6444, C => n7539, D => n7540, Z => 
                           n3998);
   U7338 : AO6 port map( A => v_RAM_IN0_11_port, B => n6538, C => n7541, Z => 
                           n7540);
   U7339 : AO4 port map( A => n7542, B => n6541, C => n7543, D => n6543, Z => 
                           n7541);
   U7340 : EO port map( A => n7544, B => n7545, Z => n7543);
   U7341 : EO port map( A => n7483, B => n7546, Z => n7545);
   U7342 : EN port map( A => n7234, B => n7231, Z => n7483);
   U7343 : EN port map( A => n4954, B => n4984, Z => n7231);
   U7344 : EN port map( A => v_KEY_COLUMN_25_port, B => n7860, Z => n4984);
   U7345 : EN port map( A => n4918, B => n4927, Z => n7234);
   U7346 : EN port map( A => v_KEY_COLUMN_9_port, B => n7868, Z => n4927);
   U7347 : EO port map( A => n7163, B => n7547, Z => n7544);
   U7348 : EN port map( A => n4863, B => n7226, Z => n7547);
   U7349 : EN port map( A => n7199, B => n4944, Z => n7226);
   U7350 : EN port map( A => v_KEY_COLUMN_18_port, B => n7931, Z => n4944);
   U7351 : EN port map( A => v_KEY_COLUMN_3_port, B => n7862, Z => n4863);
   U7352 : EO port map( A => n7548, B => n7549, Z => n7542);
   U7353 : EO port map( A => n7488, B => n7550, Z => n7549);
   U7354 : EO port map( A => n7248, B => n7244, Z => n7488);
   U7355 : EN port map( A => n5507, B => n7450, Z => n7244);
   U7356 : EO port map( A => v_KEY_COLUMN_9_port, B => n7809, Z => n7450);
   U7357 : EN port map( A => n6584, B => n7029, Z => n7248);
   U7358 : EN port map( A => v_KEY_COLUMN_25_port, B => n7936, Z => n7029);
   U7359 : EO port map( A => n7170, B => n7551, Z => n7548);
   U7360 : EN port map( A => n5257, B => n7241, Z => n7551);
   U7361 : EO port map( A => n5821, B => n6125, Z => n7241);
   U7362 : EN port map( A => v_KEY_COLUMN_18_port, B => n7874, Z => n6125);
   U7363 : EO port map( A => v_KEY_COLUMN_3_port, B => n4381, Z => n5257);
   U7364 : AO2 port map( A => n6440, B => n7552, C => n6551, D => n7553, Z => 
                           n7539);
   U7365 : EO port map( A => n7554, B => n7555, Z => n7553);
   U7366 : EO port map( A => n7495, B => n7556, Z => n7555);
   U7367 : EN port map( A => n7263, B => n7260, Z => n7495);
   U7368 : EN port map( A => n4712, B => n4727, Z => n7260);
   U7369 : EO port map( A => v_KEY_COLUMN_25_port, B => n4428, Z => n4727);
   U7370 : EN port map( A => n4621, B => n4652, Z => n7263);
   U7371 : IV port map( A => n7460, Z => n4652);
   U7372 : EO port map( A => v_KEY_COLUMN_9_port, B => n7866, Z => n7460);
   U7373 : EO port map( A => n7179, B => n7557, Z => n7554);
   U7374 : EN port map( A => n4598, B => n7255, Z => n7557);
   U7375 : EN port map( A => n7209, B => n4697, Z => n7255);
   U7376 : EN port map( A => v_KEY_COLUMN_18_port, B => n7927, Z => n4697);
   U7377 : EN port map( A => v_KEY_COLUMN_3_port, B => n7859, Z => n4598);
   U7378 : EO port map( A => v_KEY_COLUMN_11_port, B => v_DATA_COLUMN_11_port, 
                           Z => n7552);
   U7379 : EO port map( A => n7558, B => n7559, Z => n7538);
   U7380 : EO port map( A => n7500, B => n7560, Z => n7559);
   U7381 : EN port map( A => n7277, B => n7274, Z => n7500);
   U7382 : EN port map( A => n4838, B => n4848, Z => n7274);
   U7383 : IV port map( A => n7430, Z => n4848);
   U7384 : EO port map( A => v_KEY_COLUMN_25_port, B => n7863, Z => n7430);
   U7385 : EN port map( A => n4760, B => n4770, Z => n7277);
   U7386 : EN port map( A => v_KEY_COLUMN_9_port, B => n7838, Z => n4770);
   U7387 : EO port map( A => n7186, B => n7561, Z => n7558);
   U7388 : EN port map( A => n4745, B => n7269, Z => n7561);
   U7389 : EN port map( A => n7213, B => n4788, Z => n7269);
   U7390 : EN port map( A => v_KEY_COLUMN_18_port, B => n7872, Z => n4788);
   U7391 : EO port map( A => v_KEY_COLUMN_3_port, B => n4380, Z => n4745);
   U7392 : MUX21H port map( A => t_STATE_RAM0_0_11_port, B => v_RAM_IN0_11_port
                           , S => n6480, Z => n3997);
   U7393 : MUX21H port map( A => t_STATE_RAM0_1_11_port, B => v_RAM_IN0_11_port
                           , S => n6481, Z => n3996);
   U7394 : MUX21H port map( A => t_STATE_RAM0_2_11_port, B => v_RAM_IN0_11_port
                           , S => n6482, Z => n3995);
   U7395 : MUX21H port map( A => t_STATE_RAM0_3_11_port, B => v_RAM_IN0_11_port
                           , S => n4498, Z => n3994);
   U7396 : AO3 port map( A => n6483, B => n4458, C => n7562, D => n7563, Z => 
                           n3993);
   U7397 : AO2 port map( A => t_STATE_RAM0_3_11_port, B => n6486, C => 
                           v_RAM_OUT0_11_port, D => n4513, Z => n7563);
   U7398 : AO2 port map( A => t_STATE_RAM0_1_11_port, B => n4564, C => 
                           t_STATE_RAM0_2_11_port, D => n4563, Z => n7562);
   U7399 : AO3 port map( A => n7564, B => n6444, C => n7565, D => n7566, Z => 
                           n3992);
   U7400 : AO6 port map( A => v_RAM_IN0_3_port, B => n6538, C => n7567, Z => 
                           n7566);
   U7401 : AO4 port map( A => n7568, B => n6541, C => n7569, D => n6543, Z => 
                           n7567);
   U7402 : EO port map( A => n7570, B => n7571, Z => n7569);
   U7403 : EO port map( A => n7512, B => n7546, Z => n7571);
   U7404 : EO port map( A => n7513, B => n7572, Z => n7546);
   U7405 : EN port map( A => n4942, B => n4960, Z => n7572);
   U7406 : EN port map( A => v_KEY_COLUMN_27_port, B => n7816, Z => n4960);
   U7407 : EN port map( A => v_KEY_COLUMN_19_port, B => n7925, Z => n4942);
   U7408 : EN port map( A => n7573, B => n7574, Z => n7513);
   U7409 : EO port map( A => n7107, B => n7344, Z => n7574);
   U7410 : EN port map( A => n4950, B => n4986, Z => n7344);
   U7411 : IV port map( A => n7198, Z => n4950);
   U7412 : EN port map( A => n6635, B => n4929, Z => n7107);
   U7413 : EO port map( A => n6479, B => n7575, Z => n7573);
   U7414 : EO port map( A => n6478, B => n7073, Z => n7575);
   U7415 : EN port map( A => n4852, B => n7576, Z => n6479);
   U7416 : IV port map( A => n7235, Z => n4852);
   U7417 : EO port map( A => n7232, B => n7230, Z => n7512);
   U7418 : EO port map( A => n4857, B => n4888, Z => n7230);
   U7419 : EN port map( A => v_KEY_COLUMN_1_port, B => n7855, Z => n4888);
   U7420 : IV port map( A => n7381, Z => n4857);
   U7421 : EN port map( A => n6602, B => n4946, Z => n7232);
   U7422 : IV port map( A => n7443, Z => n4946);
   U7423 : EO port map( A => v_KEY_COLUMN_17_port, B => n7937, Z => n7443);
   U7424 : EO port map( A => n7163, B => n7577, Z => n7570);
   U7425 : EN port map( A => n4923, B => n7227, Z => n7577);
   U7426 : EN port map( A => n7235, B => n4865, Z => n7227);
   U7427 : EN port map( A => v_KEY_COLUMN_2_port, B => n7870, Z => n4865);
   U7428 : EN port map( A => v_KEY_COLUMN_11_port, B => n7821, Z => n4923);
   U7429 : EN port map( A => n6635, B => n4925, Z => n7163);
   U7430 : EN port map( A => v_KEY_COLUMN_10_port, B => n7820, Z => n4925);
   U7431 : IV port map( A => n6464, Z => n6541);
   U7432 : EO port map( A => n7578, B => n7579, Z => n7568);
   U7433 : EO port map( A => n7518, B => n7550, Z => n7579);
   U7434 : EO port map( A => n7519, B => n7580, Z => n7550);
   U7435 : EN port map( A => n6076, B => n6664, Z => n7580);
   U7436 : EN port map( A => v_KEY_COLUMN_27_port, B => n7924, Z => n6664);
   U7437 : EN port map( A => v_KEY_COLUMN_19_port, B => n7865, Z => n6076);
   U7438 : EN port map( A => n7581, B => n7582, Z => n7519);
   U7439 : EO port map( A => n7113, B => n7350, Z => n7582);
   U7440 : EN port map( A => n6229, B => n7307, Z => n7350);
   U7441 : EN port map( A => n5416, B => n5820, Z => n7113);
   U7442 : EO port map( A => n7082, B => n7583, Z => n7581);
   U7443 : EO port map( A => n6468, B => n7081, Z => n7583);
   U7444 : EO port map( A => n5821, B => n6199, Z => n7081);
   U7445 : EN port map( A => n5008, B => n7584, Z => n7082);
   U7446 : IV port map( A => n6472, Z => n5008);
   U7447 : EN port map( A => n7246, B => n7245, Z => n7518);
   U7448 : EN port map( A => n5095, B => n5345, Z => n7245);
   U7449 : EO port map( A => v_KEY_COLUMN_1_port, B => n4383, Z => n5345);
   U7450 : IV port map( A => n7585, Z => n5095);
   U7451 : EN port map( A => n6607, B => n6164, Z => n7246);
   U7452 : EN port map( A => v_KEY_COLUMN_17_port, B => n7873, Z => n6164);
   U7453 : EO port map( A => n7170, B => n7586, Z => n7578);
   U7454 : EN port map( A => n5671, B => n7240, Z => n7586);
   U7455 : EN port map( A => n6472, B => n5305, Z => n7240);
   U7456 : EN port map( A => v_KEY_COLUMN_2_port, B => n7932, Z => n5305);
   U7457 : EN port map( A => v_KEY_COLUMN_11_port, B => n7811, Z => n5671);
   U7458 : EN port map( A => n6643, B => n5713, Z => n7170);
   U7459 : EN port map( A => v_KEY_COLUMN_10_port, B => n7810, Z => n5713);
   U7460 : AO2 port map( A => n6440, B => n7587, C => n6551, D => n7588, Z => 
                           n7565);
   U7461 : EO port map( A => n7589, B => n7590, Z => n7588);
   U7462 : EO port map( A => n7526, B => n7556, Z => n7590);
   U7463 : EN port map( A => n7527, B => n7591, Z => n7556);
   U7464 : EN port map( A => n4694, B => n4721, Z => n7591);
   U7465 : EN port map( A => v_KEY_COLUMN_27_port, B => n7922, Z => n4721);
   U7466 : EN port map( A => v_KEY_COLUMN_19_port, B => n7921, Z => n4694);
   U7467 : EN port map( A => n7592, B => n7593, Z => n7527);
   U7468 : EN port map( A => n7119, B => n7459, Z => n7593);
   U7469 : EO port map( A => n4707, B => n4730, Z => n7459);
   U7470 : IV port map( A => n7208, Z => n4707);
   U7471 : EN port map( A => n6653, B => n4655, Z => n7119);
   U7472 : EO port map( A => n6453, B => n7594, Z => n7592);
   U7473 : EO port map( A => n6451, B => n7088, Z => n7594);
   U7474 : EN port map( A => n4583, B => n4612, Z => n6453);
   U7475 : IV port map( A => n7264, Z => n4583);
   U7476 : EN port map( A => n7261, B => n7259, Z => n7526);
   U7477 : EO port map( A => n7394, B => n4604, Z => n7259);
   U7478 : EN port map( A => v_KEY_COLUMN_1_port, B => n7853, Z => n4604);
   U7479 : EN port map( A => n6614, B => n4700, Z => n7261);
   U7480 : EO port map( A => v_KEY_COLUMN_17_port, B => n4427, Z => n4700);
   U7481 : EO port map( A => n7179, B => n7595, Z => n7589);
   U7482 : EN port map( A => n4628, B => n7256, Z => n7595);
   U7483 : EN port map( A => n7264, B => n4601, Z => n7256);
   U7484 : EN port map( A => v_KEY_COLUMN_2_port, B => n7867, Z => n4601);
   U7485 : EN port map( A => v_KEY_COLUMN_11_port, B => n7845, Z => n4628);
   U7486 : EN port map( A => n6653, B => n4631, Z => n7179);
   U7487 : EN port map( A => v_KEY_COLUMN_10_port, B => n7844, Z => n4631);
   U7488 : EO port map( A => v_KEY_COLUMN_3_port, B => v_DATA_COLUMN_3_port, Z 
                           => n7587);
   U7489 : EO port map( A => n7596, B => n7597, Z => n7564);
   U7490 : EO port map( A => n7532, B => n7560, Z => n7597);
   U7491 : EO port map( A => n7533, B => n7598, Z => n7560);
   U7492 : EN port map( A => n4786, B => n4844, Z => n7598);
   U7493 : EN port map( A => v_KEY_COLUMN_27_port, B => n7829, Z => n4844);
   U7494 : EN port map( A => v_KEY_COLUMN_19_port, B => n7864, Z => n4786);
   U7495 : EN port map( A => n7599, B => n7600, Z => n7533);
   U7496 : EO port map( A => n7125, B => n7364, Z => n7600);
   U7497 : EN port map( A => n4834, B => n4850, Z => n7364);
   U7498 : IV port map( A => n6457, Z => n4834);
   U7499 : EN port map( A => n6661, B => n4772, Z => n7125);
   U7500 : EO port map( A => n6456, B => n7601, Z => n7599);
   U7501 : EO port map( A => n6458, B => n7094, Z => n7601);
   U7502 : EN port map( A => n4734, B => n7602, Z => n6456);
   U7503 : IV port map( A => n7278, Z => n4734);
   U7504 : EO port map( A => n7275, B => n7273, Z => n7532);
   U7505 : EO port map( A => n4739, B => n4749, Z => n7273);
   U7506 : EN port map( A => v_KEY_COLUMN_1_port, B => n7935, Z => n4749);
   U7507 : IV port map( A => n7401, Z => n4739);
   U7508 : EN port map( A => n6619, B => n4810, Z => n7275);
   U7509 : IV port map( A => n7467, Z => n4810);
   U7510 : EO port map( A => v_KEY_COLUMN_17_port, B => n7833, Z => n7467);
   U7511 : EO port map( A => n7186, B => n7603, Z => n7596);
   U7512 : EN port map( A => n4765, B => n7270, Z => n7603);
   U7513 : EN port map( A => n7278, B => n4747, Z => n7270);
   U7514 : EO port map( A => v_KEY_COLUMN_2_port, B => n4382, Z => n4747);
   U7515 : EN port map( A => v_KEY_COLUMN_11_port, B => n7840, Z => n4765);
   U7516 : EN port map( A => n6661, B => n4767, Z => n7186);
   U7517 : EN port map( A => v_KEY_COLUMN_10_port, B => n7839, Z => n4767);
   U7518 : MUX21H port map( A => t_STATE_RAM0_0_3_port, B => v_RAM_IN0_3_port, 
                           S => n6480, Z => n3991);
   U7519 : MUX21H port map( A => t_STATE_RAM0_1_3_port, B => v_RAM_IN0_3_port, 
                           S => n6481, Z => n3990);
   U7520 : MUX21H port map( A => t_STATE_RAM0_2_3_port, B => v_RAM_IN0_3_port, 
                           S => n6482, Z => n3989);
   U7521 : MUX21H port map( A => t_STATE_RAM0_3_3_port, B => v_RAM_IN0_3_port, 
                           S => n4498, Z => n3988);
   U7522 : AO3 port map( A => n6483, B => n4459, C => n7604, D => n7605, Z => 
                           n3987);
   U7523 : AO2 port map( A => t_STATE_RAM0_3_3_port, B => n6486, C => 
                           v_RAM_OUT0_3_port, D => n4513, Z => n7605);
   U7524 : AO2 port map( A => t_STATE_RAM0_1_3_port, B => n4564, C => 
                           t_STATE_RAM0_2_3_port, D => n4563, Z => n7604);
   U7525 : ND4 port map( A => n7606, B => n7607, C => n7608, D => n7609, Z => 
                           n3986);
   U7526 : ND2 port map( A => n6440, B => n7610, Z => n7609);
   U7527 : EO port map( A => v_KEY_COLUMN_8_port, B => v_DATA_COLUMN_8_port, Z 
                           => n7610);
   U7528 : AO2 port map( A => n6551, B => n7611, C => n7612, D => n7613, Z => 
                           n7608);
   U7529 : EO port map( A => n7614, B => n7615, Z => n7613);
   U7530 : EO port map( A => n7094, B => n7616, Z => n7615);
   U7531 : EN port map( A => n7213, B => n4812, Z => n7094);
   U7532 : EN port map( A => n4754, B => n6461, Z => n7614);
   U7533 : EN port map( A => n4760, B => n4838, Z => n6461);
   U7534 : EN port map( A => v_KEY_COLUMN_30_port, B => n7831, Z => n4838);
   U7535 : EO port map( A => v_KEY_COLUMN_14_port, B => n7842, Z => n4760);
   U7536 : EO port map( A => n7617, B => n7618, Z => n7611);
   U7537 : EO port map( A => n7088, B => n7619, Z => n7618);
   U7538 : EN port map( A => n7209, B => n4703, Z => n7088);
   U7539 : EN port map( A => n4613, B => n6449, Z => n7617);
   U7540 : EN port map( A => n4621, B => n4712, Z => n6449);
   U7541 : EN port map( A => v_KEY_COLUMN_30_port, B => n7904, Z => n4712);
   U7542 : EO port map( A => v_KEY_COLUMN_14_port, B => n7847, Z => n4621);
   U7543 : MUX21L port map( A => n7620, B => n7621, S => n7622, Z => n7607);
   U7544 : EO port map( A => n7623, B => n7624, Z => n7622);
   U7545 : EN port map( A => n6199, B => n6470, Z => n7624);
   U7546 : EN port map( A => n6812, B => n5381, Z => n6470);
   U7547 : EN port map( A => n5507, B => n6584, Z => n6812);
   U7548 : EO port map( A => v_KEY_COLUMN_30_port, B => n7906, Z => n6584);
   U7549 : EN port map( A => v_KEY_COLUMN_14_port, B => n7813, Z => n5507);
   U7550 : EN port map( A => n6643, B => n5821, Z => n7623);
   U7551 : AO2 port map( A => n6462, B => n7625, C => v_RAM_IN0_8_port, D => 
                           n6538, Z => n7606);
   U7552 : EO port map( A => n7626, B => n7627, Z => n7625);
   U7553 : EO port map( A => n7073, B => n7628, Z => n7627);
   U7554 : EN port map( A => n7199, B => n4948, Z => n7073);
   U7555 : EN port map( A => n4912, B => n6477, Z => n7626);
   U7556 : EN port map( A => n4918, B => n4954, Z => n6477);
   U7557 : EN port map( A => v_KEY_COLUMN_30_port, B => n7818, Z => n4954);
   U7558 : EO port map( A => v_KEY_COLUMN_14_port, B => n7823, Z => n4918);
   U7559 : MUX21H port map( A => t_STATE_RAM0_0_8_port, B => v_RAM_IN0_8_port, 
                           S => n6480, Z => n3985);
   U7560 : MUX21H port map( A => t_STATE_RAM0_1_8_port, B => v_RAM_IN0_8_port, 
                           S => n6481, Z => n3984);
   U7561 : MUX21H port map( A => t_STATE_RAM0_2_8_port, B => v_RAM_IN0_8_port, 
                           S => n6482, Z => n3983);
   U7562 : MUX21H port map( A => t_STATE_RAM0_3_8_port, B => v_RAM_IN0_8_port, 
                           S => n4498, Z => n3982);
   U7563 : AO3 port map( A => n6483, B => n4460, C => n7629, D => n7630, Z => 
                           n3981);
   U7564 : AO2 port map( A => t_STATE_RAM0_3_8_port, B => n6486, C => 
                           v_RAM_OUT0_8_port, D => n4513, Z => n7630);
   U7565 : AO2 port map( A => t_STATE_RAM0_1_8_port, B => n4564, C => 
                           t_STATE_RAM0_2_8_port, D => n4563, Z => n7629);
   U7566 : AO3 port map( A => n7631, B => n6444, C => n7632, D => n7633, Z => 
                           n3980);
   U7567 : NR2 port map( A => n7634, B => n7635, Z => n7633);
   U7568 : AO4 port map( A => n6437, B => n4377, C => n7636, D => n6543, Z => 
                           n7635);
   U7569 : IV port map( A => n6462, Z => n6543);
   U7570 : EO port map( A => n7637, B => n7638, Z => n7636);
   U7571 : EN port map( A => n6782, B => n7628, Z => n7638);
   U7572 : EN port map( A => n4890, B => n7639, Z => n7628);
   U7573 : IV port map( A => n7576, Z => n4890);
   U7574 : EO port map( A => v_KEY_COLUMN_0_port, B => n7861, Z => n7576);
   U7575 : EN port map( A => n4929, B => n6631, Z => n7637);
   U7576 : EN port map( A => n7198, B => n4931, Z => n6631);
   U7577 : IV port map( A => n7199, Z => n4931);
   U7578 : EO port map( A => v_KEY_COLUMN_23_port, B => n7901, Z => n7199);
   U7579 : EO port map( A => v_KEY_COLUMN_31_port, B => n7819, Z => n7198);
   U7580 : MUX21L port map( A => n7640, B => n7641, S => n7642, Z => n7634);
   U7581 : EO port map( A => n7643, B => n7644, Z => n7642);
   U7582 : EO port map( A => n6639, B => n6777, Z => n7644);
   U7583 : EO port map( A => n5821, B => n6229, Z => n6639);
   U7584 : EN port map( A => v_KEY_COLUMN_31_port, B => n7900, Z => n6229);
   U7585 : EN port map( A => v_KEY_COLUMN_23_port, B => n7875, Z => n5821);
   U7586 : EN port map( A => n5381, B => n5820, Z => n7643);
   U7587 : IV port map( A => n7584, Z => n5381);
   U7588 : EO port map( A => v_KEY_COLUMN_0_port, B => n7944, Z => n7584);
   U7589 : AO2 port map( A => n6440, B => n7645, C => n6551, D => n7646, Z => 
                           n7632);
   U7590 : EO port map( A => n7647, B => n7648, Z => n7646);
   U7591 : EO port map( A => n6765, B => n7619, Z => n7648);
   U7592 : EO port map( A => n4612, B => n7649, Z => n7619);
   U7593 : EO port map( A => v_KEY_COLUMN_0_port, B => n7858, Z => n4612);
   U7594 : EN port map( A => n4655, B => n6649, Z => n7647);
   U7595 : EN port map( A => n7208, B => n4679, Z => n6649);
   U7596 : IV port map( A => n7209, Z => n4679);
   U7597 : EO port map( A => v_KEY_COLUMN_23_port, B => n7897, Z => n7209);
   U7598 : EO port map( A => v_KEY_COLUMN_31_port, B => n7898, Z => n7208);
   U7599 : EO port map( A => v_KEY_COLUMN_16_port, B => v_DATA_COLUMN_16_port, 
                           Z => n7645);
   U7600 : IV port map( A => n7612, Z => n6444);
   U7601 : EO port map( A => n7650, B => n7651, Z => n7631);
   U7602 : EN port map( A => n6770, B => n7616, Z => n7651);
   U7603 : EN port map( A => n4751, B => n7652, Z => n7616);
   U7604 : IV port map( A => n7602, Z => n4751);
   U7605 : EO port map( A => v_KEY_COLUMN_0_port, B => n7941, Z => n7602);
   U7606 : EN port map( A => n4772, B => n6657, Z => n7650);
   U7607 : EN port map( A => n6457, B => n4775, Z => n6657);
   U7608 : IV port map( A => n7213, Z => n4775);
   U7609 : EO port map( A => v_KEY_COLUMN_23_port, B => n7837, Z => n7213);
   U7610 : EO port map( A => v_KEY_COLUMN_31_port, B => n7832, Z => n6457);
   U7611 : MUX21L port map( A => n4426, B => n4377, S => n6480, Z => n3979);
   U7612 : MUX21H port map( A => t_STATE_RAM0_1_16_port, B => v_RAM_IN0_16_port
                           , S => n6481, Z => n3978);
   U7613 : MUX21H port map( A => t_STATE_RAM0_2_16_port, B => v_RAM_IN0_16_port
                           , S => n6482, Z => n3977);
   U7614 : MUX21H port map( A => t_STATE_RAM0_3_16_port, B => v_RAM_IN0_16_port
                           , S => n4498, Z => n3976);
   U7615 : AO3 port map( A => n6483, B => n4426, C => n7653, D => n7654, Z => 
                           n3975);
   U7616 : AO2 port map( A => t_STATE_RAM0_3_16_port, B => n6486, C => 
                           v_RAM_OUT0_16_port, D => n4513, Z => n7654);
   U7617 : AO2 port map( A => t_STATE_RAM0_1_16_port, B => n4564, C => 
                           t_STATE_RAM0_2_16_port, D => n4563, Z => n7653);
   U7618 : ND4 port map( A => n7655, B => n7656, C => n7657, D => n7658, Z => 
                           n3974);
   U7619 : ND2 port map( A => n7612, B => n7659, Z => n7658);
   U7620 : EO port map( A => n7660, B => n7661, Z => n7659);
   U7621 : EO port map( A => n6770, B => n7652, Z => n7661);
   U7622 : EN port map( A => n6458, B => n4850, Z => n7652);
   U7623 : EN port map( A => v_KEY_COLUMN_24_port, B => n7828, Z => n4850);
   U7624 : EN port map( A => n6617, B => n6656, Z => n6458);
   U7625 : EO port map( A => n4741, B => n4783, Z => n6656);
   U7626 : EO port map( A => v_KEY_COLUMN_21_port, B => n7835, Z => n4783);
   U7627 : EO port map( A => v_KEY_COLUMN_5_port, B => n4378, Z => n4741);
   U7628 : EO port map( A => n4761, B => n4840, Z => n6617);
   U7629 : EN port map( A => v_KEY_COLUMN_29_port, B => n7830, Z => n4840);
   U7630 : IV port map( A => n6806, Z => n4761);
   U7631 : EO port map( A => v_KEY_COLUMN_13_port, B => n7880, Z => n6806);
   U7632 : EN port map( A => n7401, B => n4779, Z => n6770);
   U7633 : IV port map( A => n6619, Z => n4779);
   U7634 : EO port map( A => v_KEY_COLUMN_22_port, B => n7836, Z => n6619);
   U7635 : EO port map( A => v_KEY_COLUMN_6_port, B => n7905, Z => n7401);
   U7636 : EO port map( A => n6460, B => n6574, Z => n7660);
   U7637 : EN port map( A => n7278, B => n4754, Z => n6574);
   U7638 : IV port map( A => n6661, Z => n4754);
   U7639 : EO port map( A => v_KEY_COLUMN_15_port, B => n7843, Z => n6661);
   U7640 : EO port map( A => v_KEY_COLUMN_7_port, B => n7899, Z => n7278);
   U7641 : EO port map( A => n4772, B => n4812, Z => n6460);
   U7642 : EN port map( A => v_KEY_COLUMN_16_port, B => n7878, Z => n4812);
   U7643 : EN port map( A => v_KEY_COLUMN_8_port, B => n7879, Z => n4772);
   U7644 : NR2 port map( A => n7662, B => n7663, Z => n7612);
   U7645 : AO2 port map( A => n6440, B => n7664, C => n6551, D => n7665, Z => 
                           n7657);
   U7646 : EO port map( A => n7666, B => n7667, Z => n7665);
   U7647 : EO port map( A => n6765, B => n7649, Z => n7667);
   U7648 : EN port map( A => n6451, B => n4730, Z => n7649);
   U7649 : EN port map( A => v_KEY_COLUMN_24_port, B => n7940, Z => n4730);
   U7650 : EN port map( A => n6612, B => n6648, Z => n6451);
   U7651 : EO port map( A => n4592, B => n4690, Z => n6648);
   U7652 : EO port map( A => v_KEY_COLUMN_21_port, B => n7909, Z => n4690);
   U7653 : EN port map( A => v_KEY_COLUMN_5_port, B => n7849, Z => n4592);
   U7654 : EO port map( A => n4622, B => n4715, Z => n6612);
   U7655 : EN port map( A => v_KEY_COLUMN_29_port, B => n7910, Z => n4715);
   U7656 : IV port map( A => n6799, Z => n4622);
   U7657 : EO port map( A => v_KEY_COLUMN_13_port, B => n7877, Z => n6799);
   U7658 : EN port map( A => n7394, B => n4684, Z => n6765);
   U7659 : IV port map( A => n6614, Z => n4684);
   U7660 : EO port map( A => v_KEY_COLUMN_22_port, B => n7903, Z => n6614);
   U7661 : EO port map( A => v_KEY_COLUMN_6_port, B => n7850, Z => n7394);
   U7662 : EO port map( A => n6452, B => n6569, Z => n7666);
   U7663 : EN port map( A => n7264, B => n4613, Z => n6569);
   U7664 : IV port map( A => n6653, Z => n4613);
   U7665 : EO port map( A => v_KEY_COLUMN_15_port, B => n7848, Z => n6653);
   U7666 : EO port map( A => v_KEY_COLUMN_7_port, B => n7851, Z => n7264);
   U7667 : EO port map( A => n4655, B => n4703, Z => n6452);
   U7668 : EN port map( A => v_KEY_COLUMN_16_port, B => n7939, Z => n4703);
   U7669 : EN port map( A => v_KEY_COLUMN_8_port, B => n7876, Z => n4655);
   U7670 : IV port map( A => n6446, Z => n6551);
   U7671 : ND2 port map( A => n7668, B => n7669, Z => n6446);
   U7672 : EO port map( A => v_KEY_COLUMN_0_port, B => v_DATA_COLUMN_0_port, Z 
                           => n7664);
   U7673 : AN3 port map( A => n4552, B => n6437, C => n7670, Z => n6440);
   U7674 : MUX31L port map( D0 => n7620, D1 => n7621, D2 => n7671, A => n7672, 
                           B => n6581, Z => n7656);
   U7675 : EN port map( A => n6472, B => n5416, Z => n6581);
   U7676 : IV port map( A => n6643, Z => n5416);
   U7677 : EO port map( A => v_KEY_COLUMN_15_port, B => n7814, Z => n6643);
   U7678 : EO port map( A => v_KEY_COLUMN_7_port, B => n7902, Z => n6472);
   U7679 : MUX21L port map( A => n7641, B => n7640, S => n7672, Z => n7671);
   U7680 : EN port map( A => n6777, B => n6469, Z => n7672);
   U7681 : EO port map( A => n5820, B => n6199, Z => n6469);
   U7682 : EN port map( A => v_KEY_COLUMN_16_port, B => n7806, Z => n6199);
   U7683 : EO port map( A => v_KEY_COLUMN_8_port, B => n7808, Z => n5820);
   U7684 : EN port map( A => n7585, B => n5907, Z => n6777);
   U7685 : IV port map( A => n6607, Z => n5907);
   U7686 : EO port map( A => v_KEY_COLUMN_22_port, B => n7889, Z => n6607);
   U7687 : EO port map( A => v_KEY_COLUMN_6_port, B => n7908, Z => n7585);
   U7688 : IV port map( A => n7641, Z => n7621);
   U7689 : ND2 port map( A => n7673, B => n6464, Z => n7641);
   U7690 : EN port map( A => n6468, B => n7674, Z => n7673);
   U7691 : IV port map( A => n7640, Z => n7620);
   U7692 : ND2 port map( A => n6464, B => n7675, Z => n7640);
   U7693 : EN port map( A => n6468, B => n7307, Z => n7675);
   U7694 : IV port map( A => n7674, Z => n7307);
   U7695 : EO port map( A => v_KEY_COLUMN_24_port, B => n7942, Z => n7674);
   U7696 : EN port map( A => n6937, B => n6605, Z => n6468);
   U7697 : IV port map( A => n6977, Z => n6605);
   U7698 : EO port map( A => n5575, B => n6383, Z => n6977);
   U7699 : EN port map( A => v_KEY_COLUMN_29_port, B => n7912, Z => n6383);
   U7700 : IV port map( A => n6816, Z => n5575);
   U7701 : EO port map( A => v_KEY_COLUMN_13_port, B => n7883, Z => n6816);
   U7702 : IV port map( A => n6638, Z => n6937);
   U7703 : EO port map( A => n5161, B => n6029, Z => n6638);
   U7704 : EO port map( A => v_KEY_COLUMN_21_port, B => n7890, Z => n6029);
   U7705 : EO port map( A => v_KEY_COLUMN_5_port, B => n4379, Z => n5161);
   U7706 : NR3 port map( A => n7676, B => n4399, C => n7662, Z => n6464);
   U7707 : AO2 port map( A => n6462, B => n7677, C => v_RAM_IN0_0_port, D => 
                           n6538, Z => n7655);
   U7708 : EO port map( A => n7678, B => n7679, Z => n7677);
   U7709 : EO port map( A => n6782, B => n7639, Z => n7679);
   U7710 : EN port map( A => n6478, B => n4986, Z => n7639);
   U7711 : EN port map( A => v_KEY_COLUMN_24_port, B => n7815, Z => n4986);
   U7712 : EN port map( A => n6600, B => n6630, Z => n6478);
   U7713 : EO port map( A => n4859, B => n4939, Z => n6630);
   U7714 : EO port map( A => v_KEY_COLUMN_21_port, B => n7913, Z => n4939);
   U7715 : EN port map( A => v_KEY_COLUMN_5_port, B => n7825, Z => n4859);
   U7716 : EO port map( A => n4919, B => n4956, Z => n6600);
   U7717 : EN port map( A => v_KEY_COLUMN_29_port, B => n7817, Z => n4956);
   U7718 : IV port map( A => n6823, Z => n4919);
   U7719 : EO port map( A => v_KEY_COLUMN_13_port, B => n7882, Z => n6823);
   U7720 : EN port map( A => n7381, B => n4935, Z => n6782);
   U7721 : IV port map( A => n6602, Z => n4935);
   U7722 : EO port map( A => v_KEY_COLUMN_22_port, B => n7907, Z => n6602);
   U7723 : EO port map( A => v_KEY_COLUMN_6_port, B => n7826, Z => n7381);
   U7724 : EO port map( A => n6475, B => n6587, Z => n7678);
   U7725 : EN port map( A => n7235, B => n4912, Z => n6587);
   U7726 : IV port map( A => n6635, Z => n4912);
   U7727 : EO port map( A => v_KEY_COLUMN_15_port, B => n7824, Z => n6635);
   U7728 : EO port map( A => v_KEY_COLUMN_7_port, B => n7827, Z => n7235);
   U7729 : EO port map( A => n4929, B => n4948, Z => n6475);
   U7730 : EN port map( A => v_KEY_COLUMN_16_port, B => n7943, Z => n4948);
   U7731 : EN port map( A => v_KEY_COLUMN_8_port, B => n7881, Z => n4929);
   U7732 : NR2 port map( A => n7662, B => v_CALCULATION_CNTR_0_port, Z => n6462
                           );
   U7733 : ND2 port map( A => n7668, B => n7680, Z => n7662);
   U7734 : NR3 port map( A => RESET_I, B => n7670, C => n6538, Z => n7668);
   U7735 : IV port map( A => n6437, Z => n6538);
   U7736 : AO7 port map( A => n7681, B => n4513, C => n4552, Z => n6437);
   U7737 : IV port map( A => RESET_I, Z => n4552);
   U7738 : AO6 port map( A => n7682, B => n4400, C => n7670, Z => n7681);
   U7739 : OR3 port map( A => n7669, B => n4519, C => n7676, Z => n7682);
   U7740 : NR3 port map( A => v_CNT4_0_port, B => v_CNT4_1_port, C => n4432, Z 
                           => n7670);
   U7741 : MUX21H port map( A => t_STATE_RAM0_0_0_port, B => v_RAM_IN0_0_port, 
                           S => n6480, Z => n3973);
   U7742 : NR2 port map( A => n7683, B => n7884, Z => n6480);
   U7743 : MUX21H port map( A => t_STATE_RAM0_1_0_port, B => v_RAM_IN0_0_port, 
                           S => n6481, Z => n3972);
   U7744 : NR2 port map( A => n4496, B => n7884, Z => n6481);
   U7745 : MUX21H port map( A => t_STATE_RAM0_2_0_port, B => v_RAM_IN0_0_port, 
                           S => n6482, Z => n3971);
   U7746 : NR2 port map( A => n7683, B => n4414, Z => n6482);
   U7747 : ND3 port map( A => CE_I, B => n4433, C => n7891, Z => n7683);
   U7748 : MUX21H port map( A => t_STATE_RAM0_3_0_port, B => v_RAM_IN0_0_port, 
                           S => n4498, Z => n3970);
   U7749 : NR2 port map( A => n4414, B => n4496, Z => n4498);
   U7750 : ND3 port map( A => n7891, B => CE_I, C => n7885, Z => n4496);
   U7751 : AO3 port map( A => n6483, B => n4461, C => n7684, D => n7685, Z => 
                           n3969);
   U7752 : AO2 port map( A => t_STATE_RAM0_3_0_port, B => n6486, C => 
                           v_RAM_OUT0_0_port, D => n4513, Z => n7685);
   U7753 : IV port map( A => CE_I, Z => n4513);
   U7754 : AN3 port map( A => n7888, B => CE_I, C => n7887, Z => n6486);
   U7755 : AO2 port map( A => t_STATE_RAM0_1_0_port, B => n4564, C => 
                           t_STATE_RAM0_2_0_port, D => n4563, Z => n7684);
   U7756 : NR2 port map( A => n4415, B => n4558, Z => n4563);
   U7757 : AN3 port map( A => CE_I, B => n4415, C => n7888, Z => n4564);
   U7758 : OR2 port map( A => n4558, B => n7887, Z => n6483);
   U7759 : ND2 port map( A => CE_I, B => n4434, Z => n4558);
   U7760 : AO3 port map( A => n4462, B => n5009, C => n7686, D => n7687, Z => 
                           n3968);
   U7761 : AO2 port map( A => n4911, B => n7848, C => n4753, D => n7851, Z => 
                           n7687);
   U7762 : MUX21L port map( A => DATA_O_7_port, B => n7688, S => n7689, Z => 
                           n7686);
   U7763 : ND4 port map( A => n7690, B => n7691, C => n7692, D => n7693, Z => 
                           n7688);
   U7764 : AO1 port map( A => n7694, B => n7837, C => n7695, D => n7696, Z => 
                           n7693);
   U7765 : AO4 port map( A => n4463, B => n7697, C => n4384, D => n7698, Z => 
                           n7696);
   U7766 : AO7 port map( A => n4464, B => n7699, C => n7700, Z => n7695);
   U7767 : AO2 port map( A => n7701, B => n7843, C => n7900, D => n4581, Z => 
                           n7700);
   U7768 : AO6 port map( A => n7702, B => n7824, C => n7703, Z => n7692);
   U7769 : AO4 port map( A => n4465, B => n7704, C => n4385, D => n7705, Z => 
                           n7703);
   U7770 : AO2 port map( A => n7706, B => n7819, C => n7707, D => n7814, Z => 
                           n7691);
   U7771 : AO2 port map( A => n7708, B => n7827, C => n7709, D => n7875, Z => 
                           n7690);
   U7772 : AO3 port map( A => n4466, B => n5009, C => n7710, D => n7711, Z => 
                           n3967);
   U7773 : AO2 port map( A => n4911, B => n7847, C => n4753, D => n7850, Z => 
                           n7711);
   U7774 : MUX21L port map( A => DATA_O_6_port, B => n7712, S => n7689, Z => 
                           n7710);
   U7775 : AO1 port map( A => n7713, B => n7714, C => n7715, D => n7716, Z => 
                           n7712);
   U7776 : AO1 port map( A => n7694, B => n7836, C => n7717, D => n7718, Z => 
                           n7716);
   U7777 : AO4 port map( A => n4467, B => n7697, C => n4386, D => n7698, Z => 
                           n7718);
   U7778 : AO7 port map( A => n4468, B => n7699, C => n7719, Z => n7717);
   U7779 : AO2 port map( A => n7701, B => n7842, C => n7906, D => n4581, Z => 
                           n7719);
   U7780 : AO6 port map( A => n7702, B => n7823, C => n7720, Z => n7715);
   U7781 : AO4 port map( A => n4469, B => n7704, C => n4387, D => n7705, Z => 
                           n7720);
   U7782 : AO2 port map( A => n7706, B => n7818, C => n7707, D => n7813, Z => 
                           n7714);
   U7783 : AO2 port map( A => n7708, B => n7826, C => n7709, D => n7889, Z => 
                           n7713);
   U7784 : AO3 port map( A => n4470, B => n5009, C => n7721, D => n7722, Z => 
                           n3966);
   U7785 : AO2 port map( A => n4911, B => n7877, C => n4753, D => n7849, Z => 
                           n7722);
   U7786 : MUX21L port map( A => DATA_O_5_port, B => n7723, S => n7689, Z => 
                           n7721);
   U7787 : ND4 port map( A => n7724, B => n7725, C => n7726, D => n7727, Z => 
                           n7723);
   U7788 : AO1 port map( A => n7694, B => n7835, C => n7728, D => n7729, Z => 
                           n7727);
   U7789 : AO4 port map( A => n4471, B => n7697, C => n4378, D => n7698, Z => 
                           n7729);
   U7790 : AO7 port map( A => n4472, B => n7699, C => n7730, Z => n7728);
   U7791 : AO2 port map( A => n7701, B => n7880, C => n7912, D => n4581, Z => 
                           n7730);
   U7792 : AO6 port map( A => n7702, B => n7882, C => n7731, Z => n7726);
   U7793 : AO4 port map( A => n4473, B => n7704, C => n4379, D => n7705, Z => 
                           n7731);
   U7794 : AO2 port map( A => n7706, B => n7817, C => n7707, D => n7883, Z => 
                           n7725);
   U7795 : AO2 port map( A => n7708, B => n7825, C => n7709, D => n7890, Z => 
                           n7724);
   U7796 : AO3 port map( A => n4474, B => n5009, C => n7732, D => n7733, Z => 
                           n3965);
   U7797 : AO2 port map( A => n4911, B => n7846, C => n4753, D => n7852, Z => 
                           n7733);
   U7798 : MUX21L port map( A => DATA_O_4_port, B => n7734, S => n7689, Z => 
                           n7732);
   U7799 : ND4 port map( A => n7735, B => n7736, C => n7737, D => n7738, Z => 
                           n7734);
   U7800 : AO1 port map( A => n7694, B => n7834, C => n7739, D => n7740, Z => 
                           n7738);
   U7801 : AO4 port map( A => n4475, B => n7697, C => n4388, D => n7698, Z => 
                           n7740);
   U7802 : AO7 port map( A => n4476, B => n7699, C => n7741, Z => n7739);
   U7803 : AO2 port map( A => n7701, B => n7841, C => n7918, D => n4581, Z => 
                           n7741);
   U7804 : AO6 port map( A => n7702, B => n7822, C => n7742, Z => n7737);
   U7805 : AO4 port map( A => n4477, B => n7704, C => n4389, D => n7705, Z => 
                           n7742);
   U7806 : AO2 port map( A => n7706, B => n7856, C => n7707, D => n7812, Z => 
                           n7736);
   U7807 : AO2 port map( A => n7708, B => n7854, C => n7709, D => n7807, Z => 
                           n7735);
   U7808 : AO3 port map( A => n4478, B => n5009, C => n7743, D => n7744, Z => 
                           n3964);
   U7809 : AO2 port map( A => n4911, B => n7845, C => n4753, D => n7859, Z => 
                           n7744);
   U7810 : MUX21L port map( A => DATA_O_3_port, B => n7745, S => n7689, Z => 
                           n7743);
   U7811 : ND4 port map( A => n7746, B => n7747, C => n7748, D => n7749, Z => 
                           n7745);
   U7812 : AO1 port map( A => n7694, B => n7864, C => n7750, D => n7751, Z => 
                           n7749);
   U7813 : AO4 port map( A => n4479, B => n7697, C => n4380, D => n7698, Z => 
                           n7751);
   U7814 : AO7 port map( A => n4480, B => n7699, C => n7752, Z => n7750);
   U7815 : AO2 port map( A => n7701, B => n7840, C => n7924, D => n4581, Z => 
                           n7752);
   U7816 : AO6 port map( A => n7702, B => n7821, C => n7753, Z => n7748);
   U7817 : AO4 port map( A => n4481, B => n7704, C => n4381, D => n7705, Z => 
                           n7753);
   U7818 : AO2 port map( A => n7706, B => n7816, C => n7707, D => n7811, Z => 
                           n7747);
   U7819 : AO2 port map( A => n7708, B => n7862, C => n7709, D => n7865, Z => 
                           n7746);
   U7820 : AO3 port map( A => n4482, B => n5009, C => n7754, D => n7755, Z => 
                           n3963);
   U7821 : AO2 port map( A => n4911, B => n7844, C => n4753, D => n7867, Z => 
                           n7755);
   U7822 : MUX21L port map( A => DATA_O_2_port, B => n7756, S => n7689, Z => 
                           n7754);
   U7823 : ND4 port map( A => n7757, B => n7758, C => n7759, D => n7760, Z => 
                           n7756);
   U7824 : AO1 port map( A => n7694, B => n7872, C => n7761, D => n7762, Z => 
                           n7760);
   U7825 : AO4 port map( A => n4483, B => n7697, C => n4382, D => n7698, Z => 
                           n7762);
   U7826 : AO7 port map( A => n4484, B => n7699, C => n7763, Z => n7761);
   U7827 : AO2 port map( A => n7701, B => n7839, C => n7930, D => n4581, Z => 
                           n7763);
   U7828 : AO6 port map( A => n7702, B => n7820, C => n7764, Z => n7759);
   U7829 : AO4 port map( A => n4485, B => n7704, C => n4390, D => n7705, Z => 
                           n7764);
   U7830 : AO2 port map( A => n7706, B => n7869, C => n7707, D => n7810, Z => 
                           n7758);
   U7831 : AO2 port map( A => n7708, B => n7870, C => n7709, D => n7874, Z => 
                           n7757);
   U7832 : AO3 port map( A => n4427, B => n5009, C => n7765, D => n7766, Z => 
                           n3962);
   U7833 : AO2 port map( A => n4911, B => n7866, C => n4753, D => n7853, Z => 
                           n7766);
   U7834 : MUX21L port map( A => DATA_O_1_port, B => n7767, S => n7689, Z => 
                           n7765);
   U7835 : ND4 port map( A => n7768, B => n7769, C => n7770, D => n7771, Z => 
                           n7767);
   U7836 : AO1 port map( A => n7694, B => n7833, C => n7772, D => n7773, Z => 
                           n7771);
   U7837 : AO4 port map( A => n4486, B => n7697, C => n4391, D => n7698, Z => 
                           n7773);
   U7838 : AO7 port map( A => n4428, B => n7699, C => n7774, Z => n7772);
   U7839 : AO2 port map( A => n7701, B => n7838, C => n7936, D => n4581, Z => 
                           n7774);
   U7840 : AO6 port map( A => n7702, B => n7868, C => n7775, Z => n7770);
   U7841 : AO4 port map( A => n4487, B => n7704, C => n4383, D => n7705, Z => 
                           n7775);
   U7842 : AO2 port map( A => n7706, B => n7860, C => n7707, D => n7809, Z => 
                           n7769);
   U7843 : AO2 port map( A => n7708, B => n7855, C => n7709, D => n7873, Z => 
                           n7768);
   U7844 : ND4 port map( A => n4488, B => n5009, C => n7776, D => n7777, Z => 
                           n3961);
   U7845 : AO2 port map( A => n4911, B => n7876, C => n4753, D => n7858, Z => 
                           n7777);
   U7846 : IV port map( A => n4735, Z => n4753);
   U7847 : ND2 port map( A => n7676, B => n7689, Z => n4735);
   U7848 : AN3 port map( A => n4519, B => n4399, C => n7689, Z => n4911);
   U7849 : MUX21L port map( A => DATA_O_0_port, B => n7778, S => n7689, Z => 
                           n7776);
   U7850 : ND4 port map( A => n7779, B => n7780, C => n7781, D => n7782, Z => 
                           n7778);
   U7851 : AO1 port map( A => n7694, B => n7878, C => n7783, D => n7784, Z => 
                           n7782);
   U7852 : AO4 port map( A => n4489, B => n7697, C => n4392, D => n7698, Z => 
                           n7784);
   U7853 : AO7 port map( A => n4490, B => n7699, C => n7785, Z => n7783);
   U7854 : AO2 port map( A => n7701, B => n7879, C => n7942, D => n4581, Z => 
                           n7785);
   U7855 : AO6 port map( A => n7702, B => n7881, C => n7786, Z => n7781);
   U7856 : AO4 port map( A => n4491, B => n7704, C => n4393, D => n7705, Z => 
                           n7786);
   U7857 : AO2 port map( A => n7706, B => n7815, C => n7707, D => n7808, Z => 
                           n7780);
   U7858 : IV port map( A => n7787, Z => n7707);
   U7859 : IV port map( A => n7788, Z => n7706);
   U7860 : AO2 port map( A => n7708, B => n7861, C => n7709, D => n7806, Z => 
                           n7779);
   U7861 : IV port map( A => n7789, Z => n7709);
   U7862 : IV port map( A => n7790, Z => n7708);
   U7863 : IV port map( A => n5384, Z => n5009);
   U7864 : AN3 port map( A => n4519, B => v_CALCULATION_CNTR_0_port, C => n7689
                           , Z => n5384);
   U7865 : NR2 port map( A => n4400, B => n7669, Z => n7689);
   U7866 : AO4 port map( A => n3813, B => n4584, C => n7791, D => n4400, Z => 
                           n3960);
   U7867 : NR4 port map( A => n7792, B => n7793, C => n7794, D => n7795, Z => 
                           n7791);
   U7868 : ND3 port map( A => n7704, B => n7663, C => n7705, Z => n7795);
   U7869 : ND2 port map( A => n4528, B => n7796, Z => n7705);
   U7870 : IV port map( A => n7676, Z => n7663);
   U7871 : AN3 port map( A => n7797, B => n4401, C => n6228, Z => n7676);
   U7872 : ND2 port map( A => n7798, B => n4528, Z => n7704);
   U7873 : ND4 port map( A => n7788, B => n7787, C => n7790, D => n7789, Z => 
                           n7794);
   U7874 : ND2 port map( A => n7798, B => n7797, Z => n7789);
   U7875 : ND2 port map( A => n7799, B => n7797, Z => n7790);
   U7876 : IV port map( A => n4536, Z => n7797);
   U7877 : ND2 port map( A => n7798, B => n7800, Z => n7787);
   U7878 : ND2 port map( A => n7801, B => n7796, Z => n7788);
   U7879 : OR4 port map( A => n7702, B => n7701, C => n4581, D => n4519, Z => 
                           n7793);
   U7880 : NR2 port map( A => n7802, B => v_CALCULATION_CNTR_2_port, Z => n4519
                           );
   U7881 : IV port map( A => n4571, Z => n4581);
   U7882 : ND2 port map( A => n7796, B => n7800, Z => n4571);
   U7883 : AN3 port map( A => n7803, B => n4533, C => v_CALCULATION_CNTR_1_port
                           , Z => n7796);
   U7884 : NR2 port map( A => n7802, B => n4526, Z => n7701);
   U7885 : AN2 port map( A => n7798, B => n7801, Z => n7702);
   U7886 : AN3 port map( A => n4533, B => n4405, C => n7803, Z => n7798);
   U7887 : NR2 port map( A => n4416, B => v_CALCULATION_CNTR_3_port, Z => n4533
                           );
   U7888 : ND4 port map( A => n7699, B => n7698, C => n7697, D => n7804, Z => 
                           n7792);
   U7889 : IV port map( A => n7694, Z => n7804);
   U7890 : NR2 port map( A => n4536, B => n7802, Z => n7694);
   U7891 : OR3 port map( A => v_CALCULATION_CNTR_1_port, B => n4565, C => n4401
                           , Z => n7802);
   U7892 : ND2 port map( A => v_CALCULATION_CNTR_2_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n4536);
   U7893 : ND2 port map( A => n7799, B => n7800, Z => n7697);
   U7894 : ND2 port map( A => n7799, B => n4528, Z => n7698);
   U7895 : NR2 port map( A => n4399, B => v_CALCULATION_CNTR_2_port, Z => n4528
                           );
   U7896 : ND2 port map( A => n7799, B => n7801, Z => n7699);
   U7897 : NR2 port map( A => v_CALCULATION_CNTR_0_port, B => 
                           v_CALCULATION_CNTR_2_port, Z => n7801);
   U7898 : NR2 port map( A => n4566, B => n4401, Z => n7799);
   U7899 : IV port map( A => n6228, Z => n4566);
   U7900 : IV port map( A => n4610, Z => n4584);
   U7901 : NR2 port map( A => n7680, B => n4400, Z => n4610);
   U7902 : IV port map( A => n7669, Z => n7680);
   U7903 : AN3 port map( A => n7800, B => n4401, C => n6228, Z => n7669);
   U7904 : NR2 port map( A => n4565, B => n4405, Z => n6228);
   U7905 : IV port map( A => n4526, Z => n7800);
   U7906 : ND2 port map( A => v_CALCULATION_CNTR_2_port, B => n4399, Z => n4526
                           );
   U7907 : AO7 port map( A => n4565, B => n7805, C => n4494, Z => N192);
   U7908 : OR3 port map( A => n4550, B => v_CNT4_0_port, C => n4370, Z => n4494
                           );
   U7909 : IV port map( A => VALID_DATA_I, Z => n4550);
   U7910 : ND2 port map( A => v_CALCULATION_CNTR_2_port, B => n4401, Z => n7805
                           );
   U7911 : ND2 port map( A => n7803, B => n4416, Z => n4565);
   U7912 : NR3 port map( A => v_CALCULATION_CNTR_7_port, B => 
                           v_CALCULATION_CNTR_6_port, C => 
                           v_CALCULATION_CNTR_5_port, Z => n7803);

end SYN_Behavioral;
